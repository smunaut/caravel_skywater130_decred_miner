* NGSPICE file created from decred_controller.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

.subckt decred_controller CLK_LED DATA_AVAILABLE[0] DATA_AVAILABLE[1] DATA_AVAILABLE[2]
+ DATA_AVAILABLE[3] DATA_AVAILABLE[4] DATA_FROM_HASH[0] DATA_FROM_HASH[1] DATA_FROM_HASH[2]
+ DATA_FROM_HASH[3] DATA_FROM_HASH[4] DATA_FROM_HASH[5] DATA_FROM_HASH[6] DATA_FROM_HASH[7]
+ DATA_TO_HASH[0] DATA_TO_HASH[1] DATA_TO_HASH[2] DATA_TO_HASH[3] DATA_TO_HASH[4]
+ DATA_TO_HASH[5] DATA_TO_HASH[6] DATA_TO_HASH[7] EXT_RESET_N_fromHost EXT_RESET_N_toClient
+ HASH_ADDR[0] HASH_ADDR[1] HASH_ADDR[2] HASH_ADDR[3] HASH_ADDR[4] HASH_ADDR[5] HASH_EN
+ HASH_LED ID_fromClient ID_toHost IRQ_OUT_fromClient IRQ_OUT_toHost M1_CLK_IN M1_CLK_SELECT
+ MACRO_RD_SELECT[0] MACRO_RD_SELECT[1] MACRO_RD_SELECT[2] MACRO_RD_SELECT[3] MACRO_RD_SELECT[4]
+ MACRO_WR_SELECT[0] MACRO_WR_SELECT[1] MACRO_WR_SELECT[2] MACRO_WR_SELECT[3] MACRO_WR_SELECT[4]
+ MISO_fromClient MISO_toHost MOSI_fromHost MOSI_toClient PLL_INPUT S1_CLK_IN S1_CLK_SELECT
+ SCLK_fromHost SCLK_toClient SCSN_fromHost SCSN_toClient SPI_CLK_RESET_N m1_clk_local
+ VPWR VGND
X_2037_ _2204_/CLK _2015_/Q VGND VGND VPWR VPWR DATA_TO_HASH[0] sky130_fd_sc_hd__dfxtp_4
X_2106_ _2124_/CLK _2106_/D VGND VGND VPWR VPWR ID_toHost sky130_fd_sc_hd__dfxtp_4
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1270_ _1269_/Y _2244_/Q _1048_/X VGND VGND VPWR VPWR _1271_/A sky130_fd_sc_hd__nand3_4
XFILLER_3_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1606_ _1606_/A VGND VGND VPWR VPWR _2188_/D sky130_fd_sc_hd__inv_2
XFILLER_8_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1537_ _1537_/A VGND VGND VPWR VPWR _1537_/X sky130_fd_sc_hd__buf_2
XFILLER_59_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1399_ _2138_/Q _1200_/Y _1360_/Y VGND VGND VPWR VPWR _1400_/D sky130_fd_sc_hd__or3_4
X_1468_ _1465_/Y _1972_/A _1467_/Y VGND VGND VPWR VPWR _2231_/D sky130_fd_sc_hd__a21oi_4
XFILLER_63_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1322_ _1407_/A VGND VGND VPWR VPWR _1689_/B sky130_fd_sc_hd__buf_2
X_1253_ _1248_/Y _1251_/X _1255_/A VGND VGND VPWR VPWR _1253_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_1_0_0_m1_clk_local clkbuf_0_m1_clk_local/X VGND VGND VPWR VPWR clkbuf_2_1_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1184_ _1179_/X _1180_/X _1183_/Y VGND VGND VPWR VPWR _1184_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_55_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE2_4 _1910_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1940_ _1945_/A _1940_/B _1940_/C VGND VGND VPWR VPWR _1940_/Y sky130_fd_sc_hd__nand3_4
X_1871_ _1627_/A _1871_/B VGND VGND VPWR VPWR _2137_/D sky130_fd_sc_hd__xor2_4
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1236_ _2268_/Q VGND VGND VPWR VPWR _1236_/Y sky130_fd_sc_hd__inv_2
X_1305_ _1244_/B _1068_/D _1966_/C VGND VGND VPWR VPWR _1305_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_0_m1_clk_local m1_clk_local VGND VGND VPWR VPWR clkbuf_0_m1_clk_local/X sky130_fd_sc_hd__clkbuf_16
X_1098_ _1080_/A _2262_/Q _1097_/X VGND VGND VPWR VPWR _2270_/D sky130_fd_sc_hd__o21a_4
XFILLER_52_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1167_ _1167_/A VGND VGND VPWR VPWR _1167_/X sky130_fd_sc_hd__buf_2
XFILLER_20_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2070_ _2075_/CLK _2070_/D VGND VGND VPWR VPWR _2070_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_3_3_0_m1_clk_local clkbuf_3_3_0_m1_clk_local/A VGND VGND VPWR VPWR _2061_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1021_ _2006_/Q _2008_/Q VGND VGND VPWR VPWR _1022_/A sky130_fd_sc_hd__nor2_4
X_1785_ _2139_/Q VGND VGND VPWR VPWR _1785_/Y sky130_fd_sc_hd__inv_2
X_1854_ _1854_/A _1794_/Y VGND VGND VPWR VPWR _1854_/Y sky130_fd_sc_hd__nor2_4
X_1923_ _1626_/X VGND VGND VPWR VPWR _1923_/X sky130_fd_sc_hd__buf_2
X_2199_ _2027_/CLK _1567_/X VGND VGND VPWR VPWR _2199_/Q sky130_fd_sc_hd__dfxtp_4
X_2268_ _2268_/CLK _2268_/D VGND VGND VPWR VPWR _2268_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1219_ _1209_/X _1214_/C _1202_/Y VGND VGND VPWR VPWR _1219_/X sky130_fd_sc_hd__a21o_4
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1570_ _1564_/C _1552_/A _1528_/A _2198_/Q VGND VGND VPWR VPWR _1570_/Y sky130_fd_sc_hd__nand4_4
X_2053_ _2256_/CLK _2053_/D VGND VGND VPWR VPWR _2053_/Q sky130_fd_sc_hd__dfxtp_4
X_2122_ _2130_/CLK _1908_/Y VGND VGND VPWR VPWR _2020_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1004_ _1007_/A VGND VGND VPWR VPWR _1004_/Y sky130_fd_sc_hd__inv_2
X_1768_ _1751_/X _1765_/Y _1767_/Y VGND VGND VPWR VPWR _1768_/Y sky130_fd_sc_hd__o21ai_4
X_1906_ _1176_/Y _1905_/A _1905_/Y VGND VGND VPWR VPWR _1906_/Y sky130_fd_sc_hd__o21ai_4
X_1837_ _2152_/Q _1836_/X VGND VGND VPWR VPWR _1837_/X sky130_fd_sc_hd__xor2_4
X_1699_ _1997_/A _1368_/Y _1698_/Y _1398_/X VGND VGND VPWR VPWR _1699_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_40_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1622_ _1540_/B ID_fromClient VGND VGND VPWR VPWR _1622_/X sky130_fd_sc_hd__and2_4
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1553_ _1530_/C _1552_/X _1517_/A _1542_/X _1492_/A VGND VGND VPWR VPWR _1553_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1484_ _1481_/X IRQ_OUT_fromClient VGND VGND VPWR VPWR _1484_/X sky130_fd_sc_hd__and2_4
X_2036_ _2204_/CLK _2036_/D VGND VGND VPWR VPWR _2036_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2105_ _2131_/CLK _2105_/D VGND VGND VPWR VPWR _2105_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1536_ _2202_/Q VGND VGND VPWR VPWR _1538_/B sky130_fd_sc_hd__inv_2
X_1605_ _1523_/B _1603_/Y _1604_/Y VGND VGND VPWR VPWR _1606_/A sky130_fd_sc_hd__a21o_4
X_1467_ _2175_/Q _1442_/X _1461_/X VGND VGND VPWR VPWR _1467_/Y sky130_fd_sc_hd__o21ai_4
X_1398_ _1369_/Y VGND VGND VPWR VPWR _1398_/X sky130_fd_sc_hd__buf_2
XFILLER_42_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2019_ _2187_/CLK _1910_/C VGND VGND VPWR VPWR _2019_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_12_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1321_ _1321_/A VGND VGND VPWR VPWR _1407_/A sky130_fd_sc_hd__buf_2
X_1252_ _1986_/B VGND VGND VPWR VPWR _1255_/A sky130_fd_sc_hd__inv_2
XFILLER_64_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1183_ _1152_/A _1167_/X _1560_/B VGND VGND VPWR VPWR _1183_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_3_4_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_4_9_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
X_1519_ _2195_/Q VGND VGND VPWR VPWR _1519_/Y sky130_fd_sc_hd__inv_2
XINSDIODE2_5 _1905_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1870_ _1786_/Y _1788_/Y VGND VGND VPWR VPWR _1871_/B sky130_fd_sc_hd__nor2_4
XFILLER_9_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1304_ _1300_/X _1302_/X _1303_/Y VGND VGND VPWR VPWR _1304_/Y sky130_fd_sc_hd__a21oi_4
X_1166_ _1165_/X VGND VGND VPWR VPWR _1167_/A sky130_fd_sc_hd__buf_2
X_1235_ _1186_/X _1218_/Y _1225_/Y _1232_/Y _1234_/Y VGND VGND VPWR VPWR _2249_/D
+ sky130_fd_sc_hd__a41oi_4
X_1097_ _2281_/Q _2270_/Q _1090_/X VGND VGND VPWR VPWR _1097_/X sky130_fd_sc_hd__o21a_4
X_1999_ _1598_/A _2222_/Q _1999_/C VGND VGND VPWR VPWR _1999_/Y sky130_fd_sc_hd__nor3_4
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1020_ _2006_/Q VGND VGND VPWR VPWR _1039_/A sky130_fd_sc_hd__buf_2
XFILLER_46_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1922_ _1922_/A VGND VGND VPWR VPWR _1922_/Y sky130_fd_sc_hd__inv_2
X_1853_ _1783_/B VGND VGND VPWR VPWR _1854_/A sky130_fd_sc_hd__inv_2
X_1784_ _2148_/Q _1430_/A VGND VGND VPWR VPWR _1784_/Y sky130_fd_sc_hd__nand2_4
X_2267_ _2075_/CLK _1108_/X VGND VGND VPWR VPWR _2267_/Q sky130_fd_sc_hd__dfxtp_4
X_2198_ _2027_/CLK _1572_/Y VGND VGND VPWR VPWR _2198_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_37_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1149_ _2255_/Q VGND VGND VPWR VPWR _1150_/A sky130_fd_sc_hd__buf_2
X_1218_ _1012_/Y _1158_/C _1161_/Y _1263_/A _1162_/Y VGND VGND VPWR VPWR _1218_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_20_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1003_ _1003_/A VGND VGND VPWR VPWR _1986_/D sky130_fd_sc_hd__buf_2
X_2121_ _2102_/CLK _2121_/D VGND VGND VPWR VPWR _1910_/C sky130_fd_sc_hd__dfxtp_4
X_2052_ _2163_/CLK _1681_/A VGND VGND VPWR VPWR _2047_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1905_ _1905_/A _1897_/B _1905_/C VGND VGND VPWR VPWR _1905_/Y sky130_fd_sc_hd__nand3_4
XFILLER_22_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1767_ _1767_/A _1767_/B _2036_/D VGND VGND VPWR VPWR _1767_/Y sky130_fd_sc_hd__nand3_4
XFILLER_30_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1836_ _1836_/A _2151_/Q _1838_/B _1740_/X VGND VGND VPWR VPWR _1836_/X sky130_fd_sc_hd__and4_4
X_1698_ _1679_/Y _1696_/Y _1697_/Y VGND VGND VPWR VPWR _1698_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_57_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1552_ _1552_/A _1552_/B _2199_/Q _1530_/D VGND VGND VPWR VPWR _1552_/X sky130_fd_sc_hd__and4_4
X_1621_ _1540_/B _1621_/B VGND VGND VPWR VPWR _2182_/D sky130_fd_sc_hd__and2_4
XFILLER_8_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2104_ _2131_/CLK _1946_/Y VGND VGND VPWR VPWR HASH_LED sky130_fd_sc_hd__dfxtp_4
X_1483_ _1481_/X _1483_/B VGND VGND VPWR VPWR _2225_/D sky130_fd_sc_hd__and2_4
XFILLER_62_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2035_ _2061_/CLK _2035_/D VGND VGND VPWR VPWR _2035_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_54_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1819_ _1819_/A _1825_/B _1816_/D _2158_/Q VGND VGND VPWR VPWR _1819_/Y sky130_fd_sc_hd__nand4_4
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1535_ _1532_/C VGND VGND VPWR VPWR _1539_/A sky130_fd_sc_hd__buf_2
X_1604_ _1523_/B _1603_/Y _1485_/A VGND VGND VPWR VPWR _1604_/Y sky130_fd_sc_hd__o21ai_4
X_1397_ _1357_/X _2146_/Q _1362_/X VGND VGND VPWR VPWR _1397_/Y sky130_fd_sc_hd__a21oi_4
X_1466_ _1442_/X VGND VGND VPWR VPWR _1972_/A sky130_fd_sc_hd__buf_2
X_2018_ _2256_/CLK _2018_/D VGND VGND VPWR VPWR _2018_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1320_ _1324_/A VGND VGND VPWR VPWR _1321_/A sky130_fd_sc_hd__buf_2
XFILLER_64_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1182_ _1485_/A VGND VGND VPWR VPWR _1560_/B sky130_fd_sc_hd__buf_2
X_1251_ _1264_/A VGND VGND VPWR VPWR _1251_/X sky130_fd_sc_hd__buf_2
XFILLER_64_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1518_ _2194_/Q VGND VGND VPWR VPWR _1550_/A sky130_fd_sc_hd__inv_2
X_1449_ _1438_/B _1444_/X _1309_/X VGND VGND VPWR VPWR _1449_/Y sky130_fd_sc_hd__o21ai_4
XINSDIODE2_6 _2166_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1303_ _1068_/C _1264_/X _1266_/X VGND VGND VPWR VPWR _1303_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1096_ _1080_/A _2263_/Q _1095_/X VGND VGND VPWR VPWR _1096_/X sky130_fd_sc_hd__o21a_4
XFILLER_49_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1234_ _1918_/D _1178_/X _1084_/X VGND VGND VPWR VPWR _1234_/Y sky130_fd_sc_hd__o21ai_4
X_1165_ _1249_/A _1163_/Y _1249_/C VGND VGND VPWR VPWR _1165_/X sky130_fd_sc_hd__and3_4
XFILLER_20_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1998_ _2067_/Q _2068_/Q _1998_/C VGND VGND VPWR VPWR IRQ_OUT_toHost sky130_fd_sc_hd__or3_4
XFILLER_28_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1921_ _1918_/Y _1954_/B _2116_/Q _1349_/X _1920_/Y VGND VGND VPWR VPWR _1921_/X
+ sky130_fd_sc_hd__a32o_4
X_1852_ _1852_/A _1851_/Y VGND VGND VPWR VPWR _1852_/X sky130_fd_sc_hd__xor2_4
X_1783_ _2146_/Q _1783_/B VGND VGND VPWR VPWR _1846_/A sky130_fd_sc_hd__nand2_4
X_2266_ _2075_/CLK _2266_/D VGND VGND VPWR VPWR _2266_/Q sky130_fd_sc_hd__dfxtp_4
X_2197_ _2027_/CLK _2197_/D VGND VGND VPWR VPWR _1528_/A sky130_fd_sc_hd__dfxtp_4
X_1079_ _2281_/Q VGND VGND VPWR VPWR _1080_/A sky130_fd_sc_hd__inv_2
XFILLER_40_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1148_ _1003_/A _1147_/X _2275_/Q VGND VGND VPWR VPWR _1148_/X sky130_fd_sc_hd__o21a_4
X_1217_ _1217_/A VGND VGND VPWR VPWR _1263_/A sky130_fd_sc_hd__buf_2
XFILLER_25_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2120_ _2131_/CLK _2120_/D VGND VGND VPWR VPWR _2018_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_34_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1002_ _2009_/Q VGND VGND VPWR VPWR _1003_/A sky130_fd_sc_hd__buf_2
X_2051_ _2163_/CLK _1703_/A VGND VGND VPWR VPWR _2051_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_30_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1904_ _1903_/Y VGND VGND VPWR VPWR _1905_/A sky130_fd_sc_hd__buf_2
X_1835_ _1835_/A _1834_/Y VGND VGND VPWR VPWR _1835_/X sky130_fd_sc_hd__xor2_4
X_1766_ _1607_/A VGND VGND VPWR VPWR _1767_/B sky130_fd_sc_hd__buf_2
X_1697_ _1361_/Y _2135_/Q _1371_/X VGND VGND VPWR VPWR _1697_/Y sky130_fd_sc_hd__a21oi_4
X_2249_ _2101_/CLK _2249_/D VGND VGND VPWR VPWR _2249_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1551_ _1551_/A _1519_/Y _1551_/C VGND VGND VPWR VPWR _1552_/A sky130_fd_sc_hd__nor3_4
X_1620_ _1620_/A _1610_/X VGND VGND VPWR VPWR _1620_/Y sky130_fd_sc_hd__nor2_4
X_1482_ _1481_/X _2216_/Q VGND VGND VPWR VPWR _2226_/D sky130_fd_sc_hd__and2_4
XFILLER_39_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2103_ _2101_/CLK _2103_/D VGND VGND VPWR VPWR _2103_/Q sky130_fd_sc_hd__dfxtp_4
X_2034_ _2256_/CLK _2167_/Q VGND VGND VPWR VPWR _2034_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_50_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1818_ _1812_/B _1812_/C VGND VGND VPWR VPWR _1825_/B sky130_fd_sc_hd__nor2_4
X_1749_ _1229_/X _1952_/C _1197_/X _1749_/D VGND VGND VPWR VPWR _1749_/X sky130_fd_sc_hd__and4_4
XFILLER_38_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_4_0_addressalyzerBlock.SPI_CLK clkbuf_4_5_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2130_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_42_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1534_ _1532_/Y _1533_/Y VGND VGND VPWR VPWR _1540_/A sky130_fd_sc_hd__nand2_4
X_1603_ _1602_/Y _1584_/X VGND VGND VPWR VPWR _1603_/Y sky130_fd_sc_hd__nor2_4
X_1465_ _1125_/X _1459_/A _1464_/X VGND VGND VPWR VPWR _1465_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_27_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2017_ _2187_/CLK _1913_/C VGND VGND VPWR VPWR _2017_/Q sky130_fd_sc_hd__dfxtp_4
X_1396_ _1381_/Y _1395_/Y _1358_/Y VGND VGND VPWR VPWR _1396_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_50_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1181_ _1308_/A VGND VGND VPWR VPWR _1485_/A sky130_fd_sc_hd__buf_2
X_1250_ _1249_/X VGND VGND VPWR VPWR _1264_/A sky130_fd_sc_hd__buf_2
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1517_ _1517_/A VGND VGND VPWR VPWR _1531_/A sky130_fd_sc_hd__inv_2
X_1448_ _1138_/X _2234_/Q _1447_/X VGND VGND VPWR VPWR _1448_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_55_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1379_ _1375_/X _1378_/Y VGND VGND VPWR VPWR _2239_/D sky130_fd_sc_hd__nand2_4
XFILLER_23_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1302_ _1301_/Y _1263_/X _1251_/X VGND VGND VPWR VPWR _1302_/X sky130_fd_sc_hd__o21a_4
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1233_ _1198_/X VGND VGND VPWR VPWR _1918_/D sky130_fd_sc_hd__buf_2
XFILLER_52_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1095_ _1081_/X _2271_/Q _1090_/X VGND VGND VPWR VPWR _1095_/X sky130_fd_sc_hd__o21a_4
XFILLER_37_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1164_ _1012_/Y _1213_/A _1161_/Y _1217_/A VGND VGND VPWR VPWR _1249_/C sky130_fd_sc_hd__nand4_4
XFILLER_60_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1997_ _1997_/A _2070_/Q _1997_/C _2225_/Q VGND VGND VPWR VPWR _1998_/C sky130_fd_sc_hd__or4_4
XFILLER_20_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_addressalyzerBlock.SPI_CLK clkbuf_0_addressalyzerBlock.SPI_CLK/X VGND
+ VGND VPWR VPWR clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_61_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1920_ _1920_/A VGND VGND VPWR VPWR _1920_/Y sky130_fd_sc_hd__inv_2
X_1851_ _1863_/B _1857_/D _1793_/Y _1851_/D VGND VGND VPWR VPWR _1851_/Y sky130_fd_sc_hd__nand4_4
X_1782_ _1782_/A VGND VGND VPWR VPWR _1812_/B sky130_fd_sc_hd__inv_2
X_2265_ _2075_/CLK _1112_/X VGND VGND VPWR VPWR _2265_/Q sky130_fd_sc_hd__dfxtp_4
X_2196_ _2204_/CLK _1578_/Y VGND VGND VPWR VPWR _1552_/B sky130_fd_sc_hd__dfxtp_4
X_1216_ _1205_/X _1215_/Y _1033_/X VGND VGND VPWR VPWR _2251_/D sky130_fd_sc_hd__a21oi_4
XFILLER_52_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1078_ _1620_/A _1078_/B VGND VGND VPWR VPWR _2276_/D sky130_fd_sc_hd__nor2_4
X_1147_ _1147_/A VGND VGND VPWR VPWR _1147_/X sky130_fd_sc_hd__buf_2
XFILLER_25_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2050_ _2133_/CLK _2109_/Q VGND VGND VPWR VPWR _2050_/Q sky130_fd_sc_hd__dfxtp_4
X_1001_ _2008_/Q VGND VGND VPWR VPWR _1005_/A sky130_fd_sc_hd__buf_2
X_1765_ _1772_/A _1772_/B _2272_/Q VGND VGND VPWR VPWR _1765_/Y sky130_fd_sc_hd__nand3_4
XFILLER_30_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1903_ _1902_/X VGND VGND VPWR VPWR _1903_/Y sky130_fd_sc_hd__inv_2
X_1834_ _1838_/A _1832_/C VGND VGND VPWR VPWR _1834_/Y sky130_fd_sc_hd__nand2_4
X_1696_ _1692_/X _1694_/Y _1695_/X VGND VGND VPWR VPWR _1696_/Y sky130_fd_sc_hd__a21oi_4
X_2179_ _2101_/CLK _2179_/D VGND VGND VPWR VPWR _1415_/A sky130_fd_sc_hd__dfxtp_4
X_2248_ _2101_/CLK _1241_/Y VGND VGND VPWR VPWR _2248_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1550_ _1550_/A VGND VGND VPWR VPWR _1551_/A sky130_fd_sc_hd__buf_2
X_1481_ _1772_/A VGND VGND VPWR VPWR _1481_/X sky130_fd_sc_hd__buf_2
XFILLER_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2102_ _2102_/CLK _2102_/D VGND VGND VPWR VPWR _1949_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2033_ _2028_/CLK _2166_/Q VGND VGND VPWR VPWR _2028_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_62_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1748_ _1746_/X _1747_/A _1747_/Y VGND VGND VPWR VPWR _2173_/D sky130_fd_sc_hd__a21oi_4
X_1817_ _1394_/B _1816_/Y VGND VGND VPWR VPWR _1817_/Y sky130_fd_sc_hd__xnor2_4
X_1679_ _1952_/D _1857_/A _1651_/A _1632_/X _1674_/B VGND VGND VPWR VPWR _1679_/Y
+ sky130_fd_sc_hd__o41ai_4
XFILLER_53_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1602_ _1602_/A VGND VGND VPWR VPWR _1602_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1533_ CLK_LED VGND VGND VPWR VPWR _1533_/Y sky130_fd_sc_hd__inv_2
X_1464_ _2230_/Q _1137_/A VGND VGND VPWR VPWR _1464_/X sky130_fd_sc_hd__or2_4
X_1395_ _1393_/Y _1394_/Y _1647_/A VGND VGND VPWR VPWR _1395_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_35_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2016_ _2163_/CLK _2118_/Q VGND VGND VPWR VPWR _2038_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_50_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1180_ _1291_/D _1152_/Y _1171_/Y VGND VGND VPWR VPWR _1180_/X sky130_fd_sc_hd__a21o_4
X_1516_ _1144_/Y SPI_CLK_RESET_N _1516_/C VGND VGND VPWR VPWR _2206_/D sky130_fd_sc_hd__nand3_4
X_1378_ _1377_/X _1378_/B VGND VGND VPWR VPWR _1378_/Y sky130_fd_sc_hd__nand2_4
X_1447_ _1127_/X _1447_/B VGND VGND VPWR VPWR _1447_/X sky130_fd_sc_hd__or2_4
XFILLER_55_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2281_ _2214_/CLK _1999_/Y VGND VGND VPWR VPWR _2281_/Q sky130_fd_sc_hd__dfxtp_4
X_1301_ _2269_/Q VGND VGND VPWR VPWR _1301_/Y sky130_fd_sc_hd__inv_2
X_1232_ _1227_/Y _1370_/B _1248_/B VGND VGND VPWR VPWR _1232_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_64_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1094_ _1080_/X _2264_/Q _1093_/X VGND VGND VPWR VPWR _2272_/D sky130_fd_sc_hd__o21a_4
XFILLER_37_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1163_ _1162_/Y VGND VGND VPWR VPWR _1163_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1996_ _2276_/Q MISO_fromClient _1995_/X VGND VGND VPWR VPWR MISO_toHost sky130_fd_sc_hd__o21a_4
XFILLER_9_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1850_ _1850_/A VGND VGND VPWR VPWR _1863_/B sky130_fd_sc_hd__buf_2
X_1781_ _2158_/Q VGND VGND VPWR VPWR _1781_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1146_ _2256_/Q _1506_/B _2208_/Q _1507_/A _1145_/Y VGND VGND VPWR VPWR _1146_/Y
+ sky130_fd_sc_hd__o41ai_4
X_2264_ _2075_/CLK _1114_/X VGND VGND VPWR VPWR _2264_/Q sky130_fd_sc_hd__dfxtp_4
X_2195_ _2027_/CLK _1581_/Y VGND VGND VPWR VPWR _2195_/Q sky130_fd_sc_hd__dfxtp_4
X_1215_ _1206_/X _1214_/Y _1167_/X VGND VGND VPWR VPWR _1215_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_52_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1077_ _1069_/A _1995_/B _1069_/Y _1066_/Y VGND VGND VPWR VPWR _1078_/B sky130_fd_sc_hd__o22a_4
XFILLER_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1979_ _1074_/X _1986_/C _2221_/Q _1013_/Y _1978_/Y VGND VGND VPWR VPWR _2007_/D
+ sky130_fd_sc_hd__o41ai_4
XFILLER_20_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1000_ _1069_/A VGND VGND VPWR VPWR _1071_/A sky130_fd_sc_hd__inv_2
X_1902_ _1227_/Y _1922_/A _1879_/D VGND VGND VPWR VPWR _1902_/X sky130_fd_sc_hd__and3_4
XFILLER_15_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1764_ _1751_/X _1761_/Y _1763_/Y VGND VGND VPWR VPWR _1764_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_30_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1833_ _1381_/A _1833_/B VGND VGND VPWR VPWR _2154_/D sky130_fd_sc_hd__xor2_4
XFILLER_57_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1695_ _1657_/X _2151_/Q _1356_/Y VGND VGND VPWR VPWR _1695_/X sky130_fd_sc_hd__a21o_4
X_2247_ _2247_/CLK _1260_/Y VGND VGND VPWR VPWR _1986_/B sky130_fd_sc_hd__dfxtp_4
X_2178_ _2124_/CLK _2178_/D VGND VGND VPWR VPWR _1324_/A sky130_fd_sc_hd__dfxtp_4
X_1129_ _1074_/A _2222_/Q VGND VGND VPWR VPWR _1129_/Y sky130_fd_sc_hd__nor2_4
XFILLER_25_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9_0_addressalyzerBlock.SPI_CLK clkbuf_4_9_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2250_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1480_ _1308_/A VGND VGND VPWR VPWR _1772_/A sky130_fd_sc_hd__buf_2
X_2032_ _2204_/CLK _2032_/D VGND VGND VPWR VPWR _2032_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_47_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2101_ _2101_/CLK _2101_/D VGND VGND VPWR VPWR _1726_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1678_ _1377_/X _1676_/Y _1677_/Y VGND VGND VPWR VPWR _2176_/D sky130_fd_sc_hd__o21ai_4
X_1747_ _1747_/A _1473_/A VGND VGND VPWR VPWR _1747_/Y sky130_fd_sc_hd__nor2_4
X_1816_ _1805_/B _1816_/B _1809_/C _1816_/D VGND VGND VPWR VPWR _1816_/Y sky130_fd_sc_hd__nand4_4
XFILLER_53_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1532_ _2202_/Q _1543_/A _1532_/C _2204_/Q VGND VGND VPWR VPWR _1532_/Y sky130_fd_sc_hd__nand4_4
X_1601_ _1601_/A VGND VGND VPWR VPWR _2189_/D sky130_fd_sc_hd__inv_2
XFILLER_8_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1463_ _1460_/Y _1443_/X _1462_/Y VGND VGND VPWR VPWR _2232_/D sky130_fd_sc_hd__a21oi_4
X_1394_ _1346_/X _1394_/B _1349_/X VGND VGND VPWR VPWR _1394_/Y sky130_fd_sc_hd__nand3_4
X_2015_ _2061_/CLK _2015_/D VGND VGND VPWR VPWR _2015_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_27_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_1_0_m1_clk_local clkbuf_2_1_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_3_3_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_0_0_addressalyzerBlock.SPI_CLK clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_3_1_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1515_ _1514_/Y VGND VGND VPWR VPWR _2207_/D sky130_fd_sc_hd__inv_2
X_1446_ _1441_/Y _1443_/X _1445_/Y VGND VGND VPWR VPWR _2236_/D sky130_fd_sc_hd__a21oi_4
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1377_ _1722_/A VGND VGND VPWR VPWR _1377_/X sky130_fd_sc_hd__buf_2
XFILLER_11_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1300_ _1054_/Y _1299_/Y _1292_/X VGND VGND VPWR VPWR _1300_/X sky130_fd_sc_hd__a21o_4
X_2280_ _2247_/CLK _1018_/Y VGND VGND VPWR VPWR _1069_/A sky130_fd_sc_hd__dfxtp_4
X_1231_ _1255_/D VGND VGND VPWR VPWR _1248_/B sky130_fd_sc_hd__buf_2
X_1162_ _1007_/A _1161_/Y VGND VGND VPWR VPWR _1162_/Y sky130_fd_sc_hd__nor2_4
XFILLER_64_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1093_ _1081_/X _2272_/Q _1090_/X VGND VGND VPWR VPWR _1093_/X sky130_fd_sc_hd__o21a_4
XFILLER_52_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1995_ _2223_/Q _1995_/B VGND VGND VPWR VPWR _1995_/X sky130_fd_sc_hd__or2_4
X_1429_ _1427_/Y _1428_/Y _1647_/A VGND VGND VPWR VPWR _1429_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_28_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1780_ _1754_/X _1932_/A _1779_/Y VGND VGND VPWR VPWR _1780_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2263_ _2262_/CLK _2263_/D VGND VGND VPWR VPWR _2263_/Q sky130_fd_sc_hd__dfxtp_4
X_1145_ _1144_/Y _2256_/Q SPI_CLK_RESET_N VGND VGND VPWR VPWR _1145_/Y sky130_fd_sc_hd__a21boi_4
X_2194_ _2204_/CLK _2194_/D VGND VGND VPWR VPWR _2194_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_37_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1214_ _1203_/X _1209_/X _1214_/C _1966_/C VGND VGND VPWR VPWR _1214_/Y sky130_fd_sc_hd__nor4_4
X_1076_ _2276_/Q VGND VGND VPWR VPWR _1995_/B sky130_fd_sc_hd__inv_2
X_1978_ _1769_/A _1255_/A _1474_/A _1986_/D VGND VGND VPWR VPWR _1978_/Y sky130_fd_sc_hd__nand4_4
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1901_ _1015_/A _1901_/B VGND VGND VPWR VPWR _1922_/A sky130_fd_sc_hd__nor2_4
X_1832_ _1838_/A _1798_/B _1832_/C VGND VGND VPWR VPWR _1833_/B sky130_fd_sc_hd__nand3_4
XFILLER_15_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1763_ _1767_/A _1607_/X _2170_/Q VGND VGND VPWR VPWR _1763_/Y sky130_fd_sc_hd__nand3_4
X_1694_ _1426_/A _1803_/A _1657_/X VGND VGND VPWR VPWR _1694_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_57_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2246_ _2214_/CLK _2246_/D VGND VGND VPWR VPWR _1246_/A sky130_fd_sc_hd__dfxtp_4
X_1059_ _1057_/Y _2097_/Q _1058_/Y _2095_/Q VGND VGND VPWR VPWR _1059_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_40_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1128_ _2259_/Q _1127_/X _1126_/B _1128_/D VGND VGND VPWR VPWR _1999_/C sky130_fd_sc_hd__nand4_4
X_2177_ _2176_/CLK _1656_/Y VGND VGND VPWR VPWR _1655_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_15_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_14_0_addressalyzerBlock.SPI_CLK clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2247_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_21_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2100_ _2268_/CLK _1955_/Y VGND VGND VPWR VPWR _1954_/C sky130_fd_sc_hd__dfxtp_4
X_2031_ _2027_/CLK _2036_/Q VGND VGND VPWR VPWR MACRO_WR_SELECT[4] sky130_fd_sc_hd__dfxtp_4
XFILLER_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1815_ _1814_/Y VGND VGND VPWR VPWR _2163_/D sky130_fd_sc_hd__inv_2
XFILLER_7_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1677_ _1722_/A _2176_/Q VGND VGND VPWR VPWR _1677_/Y sky130_fd_sc_hd__nand2_4
X_1746_ _1744_/Y _1398_/X _1745_/Y VGND VGND VPWR VPWR _1746_/X sky130_fd_sc_hd__a21o_4
XFILLER_26_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2229_ _2211_/CLK _2229_/D VGND VGND VPWR VPWR _2229_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1531_ _1531_/A _1537_/A VGND VGND VPWR VPWR _1543_/A sky130_fd_sc_hd__nor2_4
X_1600_ _1592_/B _1592_/A _1599_/Y VGND VGND VPWR VPWR _1601_/A sky130_fd_sc_hd__o21ai_4
XFILLER_4_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1462_ _2176_/Q _1442_/X _1461_/X VGND VGND VPWR VPWR _1462_/Y sky130_fd_sc_hd__o21ai_4
X_1393_ _1645_/A _1391_/Y _1392_/Y VGND VGND VPWR VPWR _1393_/Y sky130_fd_sc_hd__o21ai_4
X_2014_ _2250_/CLK _1977_/Y VGND VGND VPWR VPWR _1029_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1729_ _2015_/D VGND VGND VPWR VPWR _1729_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1514_ _1512_/Y _1513_/Y SPI_CLK_RESET_N VGND VGND VPWR VPWR _1514_/Y sky130_fd_sc_hd__nand3_4
X_1445_ _1378_/B _1444_/X _1309_/X VGND VGND VPWR VPWR _1445_/Y sky130_fd_sc_hd__o21ai_4
X_1376_ _2278_/Q VGND VGND VPWR VPWR _1722_/A sky130_fd_sc_hd__inv_2
XFILLER_23_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1092_ _1080_/X _2265_/Q _1091_/X VGND VGND VPWR VPWR _1092_/X sky130_fd_sc_hd__o21a_4
XFILLER_49_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1161_ _2009_/Q VGND VGND VPWR VPWR _1161_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1230_ _1230_/A _1229_/X VGND VGND VPWR VPWR _1370_/B sky130_fd_sc_hd__nor2_4
X_1994_ _1992_/Y S1_CLK_SELECT _1993_/Y VGND VGND VPWR VPWR _1994_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1428_ _1346_/X _1428_/B _1428_/C VGND VGND VPWR VPWR _1428_/Y sky130_fd_sc_hd__nand3_4
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1359_ _1319_/Y _1353_/Y _1358_/Y VGND VGND VPWR VPWR _1359_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_18_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2262_ _2262_/CLK _1119_/X VGND VGND VPWR VPWR _2262_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1213_ _1213_/A VGND VGND VPWR VPWR _1966_/C sky130_fd_sc_hd__buf_2
X_1144_ _1144_/A VGND VGND VPWR VPWR _1144_/Y sky130_fd_sc_hd__inv_2
X_2193_ _2027_/CLK _1589_/X VGND VGND VPWR VPWR _1526_/D sky130_fd_sc_hd__dfxtp_4
X_1075_ _1074_/X VGND VGND VPWR VPWR _1620_/A sky130_fd_sc_hd__buf_2
XFILLER_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1977_ _1977_/A VGND VGND VPWR VPWR _1977_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1900_ _1254_/Y _1319_/B _1887_/X _1335_/Y _1899_/X VGND VGND VPWR VPWR _1900_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1831_ _1828_/A _1830_/X VGND VGND VPWR VPWR _1831_/X sky130_fd_sc_hd__xor2_4
XFILLER_15_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1762_ _1751_/A VGND VGND VPWR VPWR _1767_/A sky130_fd_sc_hd__buf_2
X_1693_ _1816_/D VGND VGND VPWR VPWR _1803_/A sky130_fd_sc_hd__inv_2
X_2245_ _2268_/CLK _1277_/Y VGND VGND VPWR VPWR _2245_/Q sky130_fd_sc_hd__dfxtp_4
X_2176_ _2176_/CLK _2176_/D VGND VGND VPWR VPWR _2176_/Q sky130_fd_sc_hd__dfxtp_4
X_1058_ _2242_/Q VGND VGND VPWR VPWR _1058_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1127_ _2219_/Q VGND VGND VPWR VPWR _1127_/X sky130_fd_sc_hd__buf_2
XFILLER_21_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2030_ _2204_/CLK _2035_/Q VGND VGND VPWR VPWR MACRO_WR_SELECT[3] sky130_fd_sc_hd__dfxtp_4
XFILLER_47_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1745_ _2067_/Q _1360_/Y _1626_/X VGND VGND VPWR VPWR _1745_/Y sky130_fd_sc_hd__nor3_4
X_1814_ _1814_/A _1809_/Y VGND VGND VPWR VPWR _1814_/Y sky130_fd_sc_hd__nand2_4
XFILLER_7_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1676_ _2070_/Q _1368_/Y _1674_/Y _1675_/X VGND VGND VPWR VPWR _1676_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_38_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2228_ _2242_/CLK _1477_/Y VGND VGND VPWR VPWR _1007_/A sky130_fd_sc_hd__dfxtp_4
X_2159_ _2163_/CLK _1824_/X VGND VGND VPWR VPWR _1816_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_3_0_0_addressalyzerBlock.SPI_CLK clkbuf_3_1_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_4_1_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_13_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1530_ _2199_/Q _1530_/B _1530_/C _1530_/D VGND VGND VPWR VPWR _1537_/A sky130_fd_sc_hd__nand4_4
X_1461_ _1607_/A VGND VGND VPWR VPWR _1461_/X sky130_fd_sc_hd__buf_2
X_1392_ _1291_/A _2082_/Q _1428_/C _1346_/A VGND VGND VPWR VPWR _1392_/Y sky130_fd_sc_hd__a2bb2oi_4
XFILLER_4_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2013_ _2247_/CLK _2013_/D VGND VGND VPWR VPWR _2013_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_50_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1728_ _1726_/Y _1336_/X _1727_/Y VGND VGND VPWR VPWR _1728_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_58_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1659_ _2053_/D VGND VGND VPWR VPWR _1659_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1513_ _1506_/B _1509_/Y _1507_/A VGND VGND VPWR VPWR _1513_/Y sky130_fd_sc_hd__nand3_4
XFILLER_4_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1375_ _1359_/Y _1363_/Y _1374_/X VGND VGND VPWR VPWR _1375_/X sky130_fd_sc_hd__a21o_4
X_1444_ _1004_/Y VGND VGND VPWR VPWR _1444_/X sky130_fd_sc_hd__buf_2
XFILLER_55_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1091_ _1081_/X _2273_/Q _1090_/X VGND VGND VPWR VPWR _1091_/X sky130_fd_sc_hd__o21a_4
XFILLER_49_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1160_ _1022_/A _1217_/A _1007_/A VGND VGND VPWR VPWR _1249_/A sky130_fd_sc_hd__a21o_4
X_1993_ _2256_/Q S1_CLK_SELECT VGND VGND VPWR VPWR _1993_/Y sky130_fd_sc_hd__nor2_4
XFILLER_60_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1358_ _1357_/X VGND VGND VPWR VPWR _1358_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1427_ _1427_/A _1427_/B VGND VGND VPWR VPWR _1427_/Y sky130_fd_sc_hd__nand2_4
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1289_ _1285_/Y _1287_/X _1288_/Y VGND VGND VPWR VPWR _2243_/D sky130_fd_sc_hd__a21oi_4
XFILLER_43_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2261_ _2262_/CLK _1121_/X VGND VGND VPWR VPWR _2261_/Q sky130_fd_sc_hd__dfxtp_4
X_2192_ _2027_/CLK _1594_/X VGND VGND VPWR VPWR _1526_/C sky130_fd_sc_hd__dfxtp_4
X_1212_ _1212_/A VGND VGND VPWR VPWR _1214_/C sky130_fd_sc_hd__buf_2
X_1143_ _2208_/Q _1507_/A _1506_/B VGND VGND VPWR VPWR _1144_/A sky130_fd_sc_hd__nor3_4
XFILLER_37_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1074_ _1074_/A VGND VGND VPWR VPWR _1074_/X sky130_fd_sc_hd__buf_2
XFILLER_33_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1976_ _1248_/B _1026_/C _1016_/X _1975_/Y VGND VGND VPWR VPWR _1977_/A sky130_fd_sc_hd__a211o_4
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1761_ _1488_/A _1761_/B _2273_/Q VGND VGND VPWR VPWR _1761_/Y sky130_fd_sc_hd__nand3_4
X_1830_ _1836_/A _1832_/C _1828_/D VGND VGND VPWR VPWR _1830_/X sky130_fd_sc_hd__and3_4
X_1692_ _1687_/X _1690_/Y _1691_/X VGND VGND VPWR VPWR _1692_/X sky130_fd_sc_hd__a21o_4
X_2244_ _2262_/CLK _1283_/Y VGND VGND VPWR VPWR _2244_/Q sky130_fd_sc_hd__dfxtp_4
X_1126_ _1125_/X _1126_/B _1128_/D VGND VGND VPWR VPWR _1126_/Y sky130_fd_sc_hd__nand3_4
X_2175_ _2250_/CLK _1701_/Y VGND VGND VPWR VPWR _2175_/Q sky130_fd_sc_hd__dfxtp_4
X_1057_ _2244_/Q VGND VGND VPWR VPWR _1057_/Y sky130_fd_sc_hd__inv_2
X_1959_ _1407_/B _1957_/X _2274_/Q _1958_/X VGND VGND VPWR VPWR _1959_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_6_0_m1_clk_local clkbuf_2_3_0_m1_clk_local/X VGND VGND VPWR VPWR _2204_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1744_ _1725_/Y _1742_/Y _1743_/X VGND VGND VPWR VPWR _1744_/Y sky130_fd_sc_hd__o21ai_4
X_1813_ _1816_/B _1809_/C _1816_/D _1809_/D _1428_/B VGND VGND VPWR VPWR _1814_/A
+ sky130_fd_sc_hd__a41o_4
X_1675_ _1786_/A _1674_/B _1630_/X VGND VGND VPWR VPWR _1675_/X sky130_fd_sc_hd__o21a_4
X_1109_ _2266_/Q _1106_/X _1101_/X VGND VGND VPWR VPWR _1109_/X sky130_fd_sc_hd__o21a_4
XFILLER_26_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2227_ _2211_/CLK _2227_/D VGND VGND VPWR VPWR _1494_/C sky130_fd_sc_hd__dfxtp_4
X_2158_ _2256_/CLK _2158_/D VGND VGND VPWR VPWR _2158_/Q sky130_fd_sc_hd__dfxtp_4
X_2089_ _2211_/CLK DATA_FROM_HASH[4] VGND VGND VPWR VPWR _2089_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1391_ _1382_/Y _1383_/Y _1390_/Y VGND VGND VPWR VPWR _1391_/Y sky130_fd_sc_hd__a21oi_4
X_1460_ _1125_/X _2232_/Q _1459_/X VGND VGND VPWR VPWR _1460_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_35_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2012_ _2211_/CLK _2012_/D VGND VGND VPWR VPWR _2012_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_35_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1727_ _1331_/X _2109_/Q _1410_/A VGND VGND VPWR VPWR _1727_/Y sky130_fd_sc_hd__a21oi_4
X_1658_ _1426_/A _1819_/A _1657_/X VGND VGND VPWR VPWR _1658_/X sky130_fd_sc_hd__a21o_4
XFILLER_58_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1589_ _1588_/X _1560_/B _1561_/X VGND VGND VPWR VPWR _1589_/X sky130_fd_sc_hd__and3_4
XFILLER_26_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1512_ _1516_/C _2208_/Q _1508_/A VGND VGND VPWR VPWR _1512_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_4_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1374_ _1865_/A _1362_/X _1373_/Y VGND VGND VPWR VPWR _1374_/X sky130_fd_sc_hd__a21o_4
X_1443_ _1442_/X VGND VGND VPWR VPWR _1443_/X sky130_fd_sc_hd__buf_2
XFILLER_23_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1090_ _1101_/A VGND VGND VPWR VPWR _1090_/X sky130_fd_sc_hd__buf_2
XFILLER_45_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1992_ S1_CLK_IN VGND VGND VPWR VPWR _1992_/Y sky130_fd_sc_hd__inv_2
X_1288_ _1048_/X _1264_/X _1266_/X VGND VGND VPWR VPWR _1288_/Y sky130_fd_sc_hd__o21ai_4
X_1357_ _1356_/Y VGND VGND VPWR VPWR _1357_/X sky130_fd_sc_hd__buf_2
X_1426_ _1426_/A VGND VGND VPWR VPWR _1427_/B sky130_fd_sc_hd__inv_2
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1142_ _1516_/C VGND VGND VPWR VPWR _1506_/B sky130_fd_sc_hd__inv_2
X_2260_ _2262_/CLK _1123_/X VGND VGND VPWR VPWR _2260_/Q sky130_fd_sc_hd__dfxtp_4
X_2191_ _2027_/CLK _1596_/X VGND VGND VPWR VPWR _1526_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_37_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1211_ _1198_/X _1749_/D VGND VGND VPWR VPWR _1212_/A sky130_fd_sc_hd__nand2_4
XFILLER_60_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1073_ _1565_/A VGND VGND VPWR VPWR _1074_/A sky130_fd_sc_hd__buf_2
XFILLER_18_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1975_ _1039_/A _1029_/A _1005_/A VGND VGND VPWR VPWR _1975_/Y sky130_fd_sc_hd__nor3_4
X_1409_ _1409_/A _1173_/A VGND VGND VPWR VPWR _1409_/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_0_0_addressalyzerBlock.SPI_CLK clkbuf_4_1_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2102_/CLK sky130_fd_sc_hd__clkbuf_1
X_1760_ _1751_/X _1758_/Y _1759_/Y VGND VGND VPWR VPWR _2171_/D sky130_fd_sc_hd__o21ai_4
X_1691_ _1423_/X _1424_/X _1150_/A _2079_/Q VGND VGND VPWR VPWR _1691_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2243_ _2262_/CLK _2243_/D VGND VGND VPWR VPWR _1048_/A sky130_fd_sc_hd__dfxtp_4
X_1125_ _2219_/Q VGND VGND VPWR VPWR _1125_/X sky130_fd_sc_hd__buf_2
X_2174_ _2250_/CLK _2174_/D VGND VGND VPWR VPWR _1722_/B sky130_fd_sc_hd__dfxtp_4
X_1056_ _1054_/Y _1064_/A _2242_/Q _1055_/Y VGND VGND VPWR VPWR _1056_/Y sky130_fd_sc_hd__a22oi_4
X_1889_ _1651_/X _1758_/Y _1887_/X _1418_/B _1888_/X VGND VGND VPWR VPWR _2131_/D
+ sky130_fd_sc_hd__o32ai_4
X_1958_ _1958_/A VGND VGND VPWR VPWR _1958_/X sky130_fd_sc_hd__buf_2
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_5_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1743_ _1876_/B _1629_/A _1630_/B VGND VGND VPWR VPWR _1743_/X sky130_fd_sc_hd__o21a_4
X_1812_ _1781_/Y _1812_/B _1812_/C VGND VGND VPWR VPWR _1816_/B sky130_fd_sc_hd__nor3_4
X_1674_ _1674_/A _1674_/B _1674_/C VGND VGND VPWR VPWR _1674_/Y sky130_fd_sc_hd__nand3_4
X_2226_ _2211_/CLK _2226_/D VGND VGND VPWR VPWR _2226_/Q sky130_fd_sc_hd__dfxtp_4
X_1108_ _2266_/Q _1105_/X _1107_/X VGND VGND VPWR VPWR _1108_/X sky130_fd_sc_hd__o21a_4
XFILLER_53_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2088_ _2102_/CLK DATA_FROM_HASH[3] VGND VGND VPWR VPWR _2080_/D sky130_fd_sc_hd__dfxtp_4
X_2157_ _2256_/CLK _1826_/X VGND VGND VPWR VPWR _1782_/A sky130_fd_sc_hd__dfxtp_4
X_1039_ _1039_/A VGND VGND VPWR VPWR _1967_/A sky130_fd_sc_hd__inv_2
XFILLER_5_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1390_ _1386_/Y _1389_/Y _1327_/A VGND VGND VPWR VPWR _1390_/Y sky130_fd_sc_hd__a21oi_4
X_2011_ _2211_/CLK _1974_/X VGND VGND VPWR VPWR _2011_/Q sky130_fd_sc_hd__dfxtp_4
X_1588_ _1585_/Y _1586_/X _1587_/X _1526_/C _1526_/D VGND VGND VPWR VPWR _1588_/X
+ sky130_fd_sc_hd__a41o_4
X_1726_ _1726_/A VGND VGND VPWR VPWR _1726_/Y sky130_fd_sc_hd__inv_2
X_1657_ _1351_/Y VGND VGND VPWR VPWR _1657_/X sky130_fd_sc_hd__buf_2
X_2209_ _2256_/Q _2209_/D SPI_CLK_RESET_N VGND VGND VPWR VPWR _2210_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_53_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1511_ _1506_/Y _1508_/Y _1510_/Y VGND VGND VPWR VPWR _2208_/D sky130_fd_sc_hd__a21oi_4
X_1442_ _1004_/Y VGND VGND VPWR VPWR _1442_/X sky130_fd_sc_hd__buf_2
XFILLER_55_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1373_ _1369_/Y _1630_/B _2278_/Q VGND VGND VPWR VPWR _1373_/Y sky130_fd_sc_hd__nand3_4
XFILLER_23_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1709_ _1705_/X _1708_/X _1339_/X VGND VGND VPWR VPWR _1709_/X sky130_fd_sc_hd__a21o_4
XFILLER_2_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1991_ _1989_/Y M1_CLK_SELECT _1990_/Y VGND VGND VPWR VPWR m1_clk_local sky130_fd_sc_hd__a21oi_4
XFILLER_9_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1425_ _1423_/X _1424_/X VGND VGND VPWR VPWR _1426_/A sky130_fd_sc_hd__nor2_4
XFILLER_55_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1287_ _1286_/Y _1263_/X _1251_/X VGND VGND VPWR VPWR _1287_/X sky130_fd_sc_hd__o21a_4
XFILLER_36_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1356_ _1651_/A _1317_/Y VGND VGND VPWR VPWR _1356_/Y sky130_fd_sc_hd__nor2_4
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2190_ _2027_/CLK _1598_/Y VGND VGND VPWR VPWR _1586_/A sky130_fd_sc_hd__dfxtp_4
X_1072_ _1070_/X _1071_/Y _1033_/X VGND VGND VPWR VPWR _2277_/D sky130_fd_sc_hd__a21oi_4
X_1141_ _1138_/X _1139_/Y _1140_/Y VGND VGND VPWR VPWR _2257_/D sky130_fd_sc_hd__a21oi_4
X_1210_ _1230_/A VGND VGND VPWR VPWR _1749_/D sky130_fd_sc_hd__buf_2
XFILLER_60_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1974_ _1986_/C _2012_/Q _1497_/X _1037_/A VGND VGND VPWR VPWR _1974_/X sky130_fd_sc_hd__a211o_4
X_1408_ _2171_/Q _1405_/X _1328_/A _1407_/Y VGND VGND VPWR VPWR _1409_/A sky130_fd_sc_hd__a211o_4
XFILLER_43_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1339_ _1327_/A VGND VGND VPWR VPWR _1339_/X sky130_fd_sc_hd__buf_2
XFILLER_28_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1690_ _1688_/Y _1689_/Y _1150_/X VGND VGND VPWR VPWR _1690_/Y sky130_fd_sc_hd__a21oi_4
X_2242_ _2242_/CLK _1298_/Y VGND VGND VPWR VPWR _2242_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1055_ _2095_/Q VGND VGND VPWR VPWR _1055_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1124_ _2259_/Q VGND VGND VPWR VPWR _1124_/Y sky130_fd_sc_hd__inv_2
X_2173_ _2250_/CLK _2173_/D VGND VGND VPWR VPWR _1473_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1957_ _1957_/A VGND VGND VPWR VPWR _1957_/X sky130_fd_sc_hd__buf_2
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1888_ _1209_/X _1229_/X _1918_/C _1761_/B _1074_/A VGND VGND VPWR VPWR _1888_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1811_ _1807_/Y _1810_/Y VGND VGND VPWR VPWR _2164_/D sky130_fd_sc_hd__nor2_4
X_1742_ _1738_/Y _1739_/Y _1741_/Y VGND VGND VPWR VPWR _1742_/Y sky130_fd_sc_hd__a21oi_4
X_1673_ _1879_/D _1346_/X _1673_/C _1952_/A VGND VGND VPWR VPWR _1674_/C sky130_fd_sc_hd__nand4_4
XFILLER_38_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2225_ _2224_/CLK _2225_/D VGND VGND VPWR VPWR _2225_/Q sky130_fd_sc_hd__dfxtp_4
X_1107_ _2267_/Q _1106_/X _1101_/X VGND VGND VPWR VPWR _1107_/X sky130_fd_sc_hd__o21a_4
X_2087_ _2130_/CLK DATA_FROM_HASH[2] VGND VGND VPWR VPWR _2087_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2156_ _2163_/CLK _1829_/X VGND VGND VPWR VPWR _2156_/Q sky130_fd_sc_hd__dfxtp_4
X_1038_ _1035_/X _1038_/B VGND VGND VPWR VPWR _1038_/X sky130_fd_sc_hd__and2_4
XFILLER_44_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2010_ _2242_/CLK _2010_/D VGND VGND VPWR VPWR _1147_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_3_2_0_m1_clk_local clkbuf_3_3_0_m1_clk_local/A VGND VGND VPWR VPWR _2256_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1725_ _1936_/B _1863_/A _1651_/A _1632_/X _1629_/A VGND VGND VPWR VPWR _1725_/Y
+ sky130_fd_sc_hd__o41ai_4
X_1587_ _1526_/A VGND VGND VPWR VPWR _1587_/X sky130_fd_sc_hd__buf_2
X_1656_ _1654_/Y _1747_/A _1655_/Y VGND VGND VPWR VPWR _1656_/Y sky130_fd_sc_hd__a21oi_4
X_2208_ _2061_/CLK _2208_/D VGND VGND VPWR VPWR _2208_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_26_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2139_ _2133_/CLK _1867_/X VGND VGND VPWR VPWR _2139_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_41_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1510_ _1516_/C _1509_/Y SPI_CLK_RESET_N VGND VGND VPWR VPWR _1510_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_4_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1441_ _1138_/X _1447_/B _1440_/X VGND VGND VPWR VPWR _1441_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_48_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1372_ _1371_/X VGND VGND VPWR VPWR _1630_/B sky130_fd_sc_hd__inv_2
X_1708_ _2118_/Q _1414_/X _1415_/X _1707_/Y VGND VGND VPWR VPWR _1708_/X sky130_fd_sc_hd__a211o_4
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1639_ _1405_/X _1639_/B VGND VGND VPWR VPWR _1639_/Y sky130_fd_sc_hd__nor2_4
XFILLER_64_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1990_ PLL_INPUT M1_CLK_SELECT VGND VGND VPWR VPWR _1990_/Y sky130_fd_sc_hd__nor2_4
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1355_ _1952_/A VGND VGND VPWR VPWR _1651_/A sky130_fd_sc_hd__inv_2
X_1424_ _1367_/Y VGND VGND VPWR VPWR _1424_/X sky130_fd_sc_hd__buf_2
XFILLER_63_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1286_ _2271_/Q VGND VGND VPWR VPWR _1286_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_5_0_addressalyzerBlock.SPI_CLK clkbuf_4_5_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2073_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_49_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1071_ _1071_/A _1071_/B VGND VGND VPWR VPWR _1071_/Y sky130_fd_sc_hd__nand2_4
X_1140_ _1138_/X _1139_/Y _1129_/Y VGND VGND VPWR VPWR _1140_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1973_ _1972_/Y _1041_/B _1476_/A VGND VGND VPWR VPWR _2012_/D sky130_fd_sc_hd__a21oi_4
X_1338_ _1335_/Y _1336_/X _1337_/Y VGND VGND VPWR VPWR _1338_/Y sky130_fd_sc_hd__o21ai_4
X_1407_ _1407_/A _1407_/B VGND VGND VPWR VPWR _1407_/Y sky130_fd_sc_hd__nor2_4
XFILLER_45_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1269_ _1278_/B VGND VGND VPWR VPWR _1269_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2172_ _2130_/CLK _2172_/D VGND VGND VPWR VPWR _1755_/C sky130_fd_sc_hd__dfxtp_4
X_2241_ _2268_/CLK _1304_/Y VGND VGND VPWR VPWR _1054_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1123_ _1105_/A _2214_/Q _1122_/X VGND VGND VPWR VPWR _1123_/X sky130_fd_sc_hd__o21a_4
X_1054_ _1054_/A VGND VGND VPWR VPWR _1054_/Y sky130_fd_sc_hd__inv_2
X_1887_ _1887_/A VGND VGND VPWR VPWR _1887_/X sky130_fd_sc_hd__buf_2
X_1956_ _1229_/X _1918_/C _1757_/A _1952_/D _1565_/A VGND VGND VPWR VPWR _1957_/A
+ sky130_fd_sc_hd__a41o_4
XFILLER_21_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1741_ _1749_/D _1740_/X _1936_/B _1198_/X _1632_/X VGND VGND VPWR VPWR _1741_/Y
+ sky130_fd_sc_hd__a2111oi_4
X_1810_ _1810_/A _1809_/Y VGND VGND VPWR VPWR _1810_/Y sky130_fd_sc_hd__nor2_4
XFILLER_7_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1672_ _1658_/X _1670_/Y _1671_/X VGND VGND VPWR VPWR _1674_/A sky130_fd_sc_hd__o21ai_4
X_1106_ _1104_/A VGND VGND VPWR VPWR _1106_/X sky130_fd_sc_hd__buf_2
X_2155_ _2163_/CLK _1831_/X VGND VGND VPWR VPWR _1828_/A sky130_fd_sc_hd__dfxtp_4
X_2224_ _2224_/CLK _1484_/X VGND VGND VPWR VPWR _1483_/B sky130_fd_sc_hd__dfxtp_4
X_2086_ _2073_/CLK DATA_FROM_HASH[1] VGND VGND VPWR VPWR _2078_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_61_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1037_ _1037_/A VGND VGND VPWR VPWR _1038_/B sky130_fd_sc_hd__inv_2
X_1939_ _1939_/A VGND VGND VPWR VPWR _1945_/A sky130_fd_sc_hd__buf_2
XFILLER_21_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_addressalyzerBlock.SPI_CLK clkbuf_0_addressalyzerBlock.SPI_CLK/X VGND
+ VGND VPWR VPWR clkbuf_2_3_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_4_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1724_ _1861_/A VGND VGND VPWR VPWR _1863_/A sky130_fd_sc_hd__inv_2
X_1586_ _1586_/A VGND VGND VPWR VPWR _1586_/X sky130_fd_sc_hd__buf_2
X_1655_ _1747_/A _1655_/B VGND VGND VPWR VPWR _1655_/Y sky130_fd_sc_hd__nor2_4
X_2207_ _2061_/CLK _2207_/D VGND VGND VPWR VPWR _1507_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_26_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2138_ _2028_/CLK _1869_/X VGND VGND VPWR VPWR _2138_/Q sky130_fd_sc_hd__dfxtp_4
X_2069_ _2102_/CLK _2074_/Q VGND VGND VPWR VPWR _1997_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1440_ _1127_/X _1486_/B VGND VGND VPWR VPWR _1440_/X sky130_fd_sc_hd__or2_4
X_1371_ _1371_/A VGND VGND VPWR VPWR _1371_/X sky130_fd_sc_hd__buf_2
XFILLER_63_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1638_ _1638_/A VGND VGND VPWR VPWR _1639_/B sky130_fd_sc_hd__inv_2
X_1707_ _1418_/A _1707_/B VGND VGND VPWR VPWR _1707_/Y sky130_fd_sc_hd__nor2_4
X_1569_ _2198_/Q _1568_/X _1485_/A VGND VGND VPWR VPWR _1569_/X sky130_fd_sc_hd__o21a_4
XFILLER_22_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1285_ _1048_/X _1269_/Y _1284_/X VGND VGND VPWR VPWR _1285_/Y sky130_fd_sc_hd__o21ai_4
X_1423_ _1344_/Y VGND VGND VPWR VPWR _1423_/X sky130_fd_sc_hd__buf_2
X_1354_ _1198_/X _1230_/A VGND VGND VPWR VPWR _1952_/A sky130_fd_sc_hd__nor2_4
XFILLER_51_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_10_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2224_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_54_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1070_ _1066_/Y _1068_/Y _1069_/Y VGND VGND VPWR VPWR _1070_/X sky130_fd_sc_hd__a21o_4
XFILLER_1_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1972_ _1972_/A _2012_/Q VGND VGND VPWR VPWR _1972_/Y sky130_fd_sc_hd__nand2_4
X_1337_ _1336_/A _2132_/Q _1415_/A VGND VGND VPWR VPWR _1337_/Y sky130_fd_sc_hd__a21oi_4
X_1406_ _2099_/Q VGND VGND VPWR VPWR _1407_/B sky130_fd_sc_hd__inv_2
X_1268_ _1262_/Y _1265_/X _1267_/Y VGND VGND VPWR VPWR _2246_/D sky130_fd_sc_hd__a21oi_4
XFILLER_28_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1199_ _2248_/Q VGND VGND VPWR VPWR _1230_/A sky130_fd_sc_hd__buf_2
XFILLER_59_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1122_ _2260_/Q _1104_/A _1115_/X VGND VGND VPWR VPWR _1122_/X sky130_fd_sc_hd__o21a_4
X_2171_ _2130_/CLK _2171_/D VGND VGND VPWR VPWR _2171_/Q sky130_fd_sc_hd__dfxtp_4
X_2240_ _2268_/CLK _2240_/D VGND VGND VPWR VPWR _1244_/D sky130_fd_sc_hd__dfxtp_4
X_1053_ _1051_/Y _2096_/Q _2245_/Q _1052_/Y VGND VGND VPWR VPWR _1060_/B sky130_fd_sc_hd__a22oi_4
X_1955_ _1254_/Y _1953_/Y _1954_/Y VGND VGND VPWR VPWR _1955_/Y sky130_fd_sc_hd__o21ai_4
X_1886_ _1885_/Y VGND VGND VPWR VPWR _1887_/A sky130_fd_sc_hd__inv_2
XFILLER_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1740_ _1740_/A VGND VGND VPWR VPWR _1740_/X sky130_fd_sc_hd__buf_2
X_1671_ _1749_/D _2152_/Q _1918_/D _1318_/X VGND VGND VPWR VPWR _1671_/X sky130_fd_sc_hd__a211o_4
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1105_ _1105_/A VGND VGND VPWR VPWR _1105_/X sky130_fd_sc_hd__buf_2
XFILLER_53_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2085_ _2176_/CLK DATA_FROM_HASH[0] VGND VGND VPWR VPWR _2077_/D sky130_fd_sc_hd__dfxtp_4
X_2154_ _2163_/CLK _2154_/D VGND VGND VPWR VPWR _1798_/A sky130_fd_sc_hd__dfxtp_4
X_2223_ _2211_/CLK _1486_/X VGND VGND VPWR VPWR _2223_/Q sky130_fd_sc_hd__dfxtp_4
X_1036_ _1039_/A _2008_/Q _1026_/C VGND VGND VPWR VPWR _1037_/A sky130_fd_sc_hd__nor3_4
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1938_ _1939_/A VGND VGND VPWR VPWR _1938_/X sky130_fd_sc_hd__buf_2
X_1869_ _2138_/Q _1868_/Y VGND VGND VPWR VPWR _1869_/X sky130_fd_sc_hd__xor2_4
XFILLER_52_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1654_ _1997_/C _1626_/X _1360_/Y _1631_/Y _1653_/Y VGND VGND VPWR VPWR _1654_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1723_ _1377_/X _1721_/Y _1722_/Y VGND VGND VPWR VPWR _2174_/D sky130_fd_sc_hd__o21ai_4
XFILLER_58_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2206_ _2256_/CLK _2206_/D VGND VGND VPWR VPWR _1516_/C sky130_fd_sc_hd__dfxtp_4
X_1585_ _1525_/A _1525_/C _1584_/X VGND VGND VPWR VPWR _1585_/Y sky130_fd_sc_hd__nor3_4
X_2068_ _2075_/CLK _2068_/D VGND VGND VPWR VPWR _2068_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_26_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2137_ _2028_/CLK _2137_/D VGND VGND VPWR VPWR _1627_/A sky130_fd_sc_hd__dfxtp_4
X_1019_ _2011_/Q VGND VGND VPWR VPWR _1026_/C sky130_fd_sc_hd__inv_2
XFILLER_1_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1370_ _1366_/Y _1370_/B _1315_/Y _1344_/B VGND VGND VPWR VPWR _1371_/A sky130_fd_sc_hd__and4_4
XFILLER_63_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1706_ _2126_/Q VGND VGND VPWR VPWR _1707_/B sky130_fd_sc_hd__inv_2
X_1637_ _1637_/A VGND VGND VPWR VPWR _1637_/Y sky130_fd_sc_hd__inv_2
X_1568_ _1564_/A _1564_/B _1552_/B _1528_/A VGND VGND VPWR VPWR _1568_/X sky130_fd_sc_hd__and4_4
X_1499_ _1497_/X SCSN_fromHost VGND VGND VPWR VPWR _2217_/D sky130_fd_sc_hd__or2_4
XFILLER_54_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1422_ _1409_/Y _1420_/Y _1421_/Y VGND VGND VPWR VPWR _1427_/A sky130_fd_sc_hd__o21ai_4
X_1284_ _1051_/Y _1278_/B _1248_/B VGND VGND VPWR VPWR _1284_/X sky130_fd_sc_hd__o21a_4
X_1353_ _1348_/Y _1350_/Y _1647_/A VGND VGND VPWR VPWR _1353_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_63_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1971_ _1967_/Y _1969_/Y _1497_/X _1970_/Y VGND VGND VPWR VPWR _1971_/X sky130_fd_sc_hd__a211o_4
X_1405_ _1321_/A VGND VGND VPWR VPWR _1405_/X sky130_fd_sc_hd__buf_2
XFILLER_5_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1336_ _1336_/A VGND VGND VPWR VPWR _1336_/X sky130_fd_sc_hd__buf_2
X_1267_ _1246_/X _1257_/X _1266_/X VGND VGND VPWR VPWR _1267_/Y sky130_fd_sc_hd__o21ai_4
X_1198_ _2249_/Q VGND VGND VPWR VPWR _1198_/X sky130_fd_sc_hd__buf_2
XFILLER_61_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_addressalyzerBlock.SPI_CLK _1994_/Y VGND VGND VPWR VPWR clkbuf_0_addressalyzerBlock.SPI_CLK/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_10_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1121_ _2260_/Q _1105_/A _1120_/X VGND VGND VPWR VPWR _1121_/X sky130_fd_sc_hd__o21a_4
X_2170_ _2073_/CLK _1764_/Y VGND VGND VPWR VPWR _2170_/Q sky130_fd_sc_hd__dfxtp_4
X_1052_ _2098_/Q VGND VGND VPWR VPWR _1052_/Y sky130_fd_sc_hd__inv_2
X_1954_ _1953_/Y _1954_/B _1954_/C VGND VGND VPWR VPWR _1954_/Y sky130_fd_sc_hd__nand3_4
XFILLER_14_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_addressalyzerBlock.SPI_CLK clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
X_1885_ _1015_/A _1936_/B _1901_/B VGND VGND VPWR VPWR _1885_/Y sky130_fd_sc_hd__nor3_4
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1319_ _1319_/A _1319_/B _1318_/X VGND VGND VPWR VPWR _1319_/Y sky130_fd_sc_hd__nor3_4
XFILLER_24_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1670_ _1668_/Y _1291_/A _1669_/X VGND VGND VPWR VPWR _1670_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_7_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2222_ _2247_/CLK _2222_/D VGND VGND VPWR VPWR _2222_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1104_ _1104_/A VGND VGND VPWR VPWR _1105_/A sky130_fd_sc_hd__inv_2
X_2084_ _2102_/CLK _2084_/D VGND VGND VPWR VPWR _2084_/Q sky130_fd_sc_hd__dfxtp_4
X_2153_ _2163_/CLK _1835_/X VGND VGND VPWR VPWR _1798_/B sky130_fd_sc_hd__dfxtp_4
X_1035_ _1028_/Y _1966_/B _1031_/X VGND VGND VPWR VPWR _1035_/X sky130_fd_sc_hd__a21o_4
XFILLER_21_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1937_ _1936_/Y VGND VGND VPWR VPWR _1939_/A sky130_fd_sc_hd__inv_2
X_1799_ _1799_/A VGND VGND VPWR VPWR _1828_/D sky130_fd_sc_hd__inv_2
X_1868_ _1627_/Y _1786_/Y _1788_/Y VGND VGND VPWR VPWR _1868_/Y sky130_fd_sc_hd__nor3_4
XFILLER_29_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1584_ _1584_/A VGND VGND VPWR VPWR _1584_/X sky130_fd_sc_hd__buf_2
X_1653_ _1648_/Y _1650_/X _1652_/Y VGND VGND VPWR VPWR _1653_/Y sky130_fd_sc_hd__a21oi_4
X_1722_ _1722_/A _1722_/B VGND VGND VPWR VPWR _1722_/Y sky130_fd_sc_hd__nand2_4
X_2205_ _2204_/CLK _2205_/D VGND VGND VPWR VPWR CLK_LED sky130_fd_sc_hd__dfxtp_4
X_2067_ _2075_/CLK _2067_/D VGND VGND VPWR VPWR _2067_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1018_ _1071_/A _1010_/Y _1017_/X VGND VGND VPWR VPWR _1018_/Y sky130_fd_sc_hd__a21oi_4
X_2136_ _2028_/CLK _1872_/X VGND VGND VPWR VPWR _1786_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_43_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1705_ _1949_/C _1414_/X _1410_/X _1704_/Y VGND VGND VPWR VPWR _1705_/X sky130_fd_sc_hd__a211o_4
XFILLER_31_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1567_ _2199_/Q _1564_/X _1566_/Y VGND VGND VPWR VPWR _1567_/X sky130_fd_sc_hd__o21a_4
XFILLER_58_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1636_ _2036_/D _1635_/A _1328_/A _1635_/Y VGND VGND VPWR VPWR _1637_/A sky130_fd_sc_hd__a211o_4
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2119_ _2101_/CLK _2119_/D VGND VGND VPWR VPWR _1913_/C sky130_fd_sc_hd__dfxtp_4
X_1498_ _1497_/X _2217_/Q VGND VGND VPWR VPWR _2218_/D sky130_fd_sc_hd__or2_4
XFILLER_14_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_15_0_addressalyzerBlock.SPI_CLK clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2242_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1421_ _1150_/X _2083_/Q VGND VGND VPWR VPWR _1421_/Y sky130_fd_sc_hd__nand2_4
XFILLER_55_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1283_ _1280_/X _1281_/X _1282_/Y VGND VGND VPWR VPWR _1283_/Y sky130_fd_sc_hd__a21oi_4
X_1352_ _1351_/Y VGND VGND VPWR VPWR _1647_/A sky130_fd_sc_hd__buf_2
XFILLER_63_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1619_ _1610_/X _1611_/X _1618_/Y VGND VGND VPWR VPWR _1619_/X sky130_fd_sc_hd__o21a_4
XFILLER_42_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1970_ _2222_/Q _1012_/Y VGND VGND VPWR VPWR _1970_/Y sky130_fd_sc_hd__nor2_4
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1335_ _2022_/D VGND VGND VPWR VPWR _1335_/Y sky130_fd_sc_hd__inv_2
X_1404_ _1647_/A _1828_/A _1357_/X VGND VGND VPWR VPWR _1404_/X sky130_fd_sc_hd__a21o_4
XFILLER_56_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1266_ _1485_/A VGND VGND VPWR VPWR _1266_/X sky130_fd_sc_hd__buf_2
XFILLER_24_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1197_ _2250_/Q VGND VGND VPWR VPWR _1197_/X sky130_fd_sc_hd__buf_2
XFILLER_51_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1120_ _2261_/Q _1104_/A _1115_/X VGND VGND VPWR VPWR _1120_/X sky130_fd_sc_hd__o21a_4
X_1051_ _1048_/A VGND VGND VPWR VPWR _1051_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1884_ _1920_/A _1881_/X _1883_/Y VGND VGND VPWR VPWR _1884_/Y sky130_fd_sc_hd__o21ai_4
X_1953_ _1958_/A VGND VGND VPWR VPWR _1953_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1318_ _1317_/Y VGND VGND VPWR VPWR _1318_/X sky130_fd_sc_hd__buf_2
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1249_ _1249_/A _1161_/Y _1249_/C VGND VGND VPWR VPWR _1249_/X sky130_fd_sc_hd__and3_4
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2221_ _2247_/CLK _1493_/Y VGND VGND VPWR VPWR _2221_/Q sky130_fd_sc_hd__dfxtp_4
X_2152_ _2133_/CLK _1837_/X VGND VGND VPWR VPWR _2152_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1103_ _1080_/A _2260_/Q _1102_/X VGND VGND VPWR VPWR _2268_/D sky130_fd_sc_hd__o21a_4
XFILLER_38_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2083_ _2176_/CLK _2091_/Q VGND VGND VPWR VPWR _2083_/Q sky130_fd_sc_hd__dfxtp_4
X_1034_ _1026_/X _1032_/X _1033_/X VGND VGND VPWR VPWR _2279_/D sky130_fd_sc_hd__a21oi_4
X_1867_ _1849_/C _1843_/Y VGND VGND VPWR VPWR _1867_/X sky130_fd_sc_hd__xor2_4
XFILLER_21_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1936_ _1015_/A _1936_/B _1901_/B _1212_/A VGND VGND VPWR VPWR _1936_/Y sky130_fd_sc_hd__nor4_4
X_1798_ _1798_/A _1798_/B VGND VGND VPWR VPWR _1799_/A sky130_fd_sc_hd__nand2_4
XFILLER_52_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1721_ _2068_/Q _1368_/Y _1720_/X _1398_/X VGND VGND VPWR VPWR _1721_/Y sky130_fd_sc_hd__a22oi_4
X_1583_ _1551_/A _1561_/X _1582_/Y VGND VGND VPWR VPWR _2194_/D sky130_fd_sc_hd__a21oi_4
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1652_ _1952_/D _1783_/B _1651_/X _1632_/X _1674_/B VGND VGND VPWR VPWR _1652_/Y
+ sky130_fd_sc_hd__o41ai_4
X_2204_ _2204_/CLK _1546_/X VGND VGND VPWR VPWR _2204_/Q sky130_fd_sc_hd__dfxtp_4
X_2135_ _2133_/CLK _1875_/Y VGND VGND VPWR VPWR _2135_/Q sky130_fd_sc_hd__dfxtp_4
X_2066_ _2061_/CLK _2066_/D VGND VGND VPWR VPWR _2066_/Q sky130_fd_sc_hd__dfxtp_4
X_1017_ _1009_/Y _1014_/Y _1016_/X VGND VGND VPWR VPWR _1017_/X sky130_fd_sc_hd__a21o_4
XFILLER_22_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1919_ _1488_/A VGND VGND VPWR VPWR _1954_/B sky130_fd_sc_hd__buf_2
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1704_ _1418_/A _1704_/B VGND VGND VPWR VPWR _1704_/Y sky130_fd_sc_hd__nor2_4
X_1566_ _1564_/C _1552_/A _2199_/Q _1530_/D _1565_/X VGND VGND VPWR VPWR _1566_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_58_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1635_ _1635_/A _1047_/Y VGND VGND VPWR VPWR _1635_/Y sky130_fd_sc_hd__nor2_4
X_1497_ _1492_/A VGND VGND VPWR VPWR _1497_/X sky130_fd_sc_hd__buf_2
X_2118_ _2102_/CLK _2118_/D VGND VGND VPWR VPWR _2118_/Q sky130_fd_sc_hd__dfxtp_4
X_2049_ _2163_/CLK _2049_/D VGND VGND VPWR VPWR MACRO_RD_SELECT[4] sky130_fd_sc_hd__dfxtp_4
XFILLER_13_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1420_ _1413_/X _1419_/X _1339_/X VGND VGND VPWR VPWR _1420_/Y sky130_fd_sc_hd__a21oi_4
X_1351_ _1313_/Y _1317_/Y VGND VGND VPWR VPWR _1351_/Y sky130_fd_sc_hd__nor2_4
XFILLER_63_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1282_ _2244_/Q _1257_/X _1266_/X VGND VGND VPWR VPWR _1282_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_36_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1618_ _1610_/X _1611_/X _1074_/X VGND VGND VPWR VPWR _1618_/Y sky130_fd_sc_hd__a21oi_4
X_1549_ _1539_/A _1539_/B _1548_/Y VGND VGND VPWR VPWR _2203_/D sky130_fd_sc_hd__o21a_4
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_1_0_addressalyzerBlock.SPI_CLK clkbuf_3_1_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_4_3_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1265_ _1176_/Y _1263_/X _1264_/X VGND VGND VPWR VPWR _1265_/X sky130_fd_sc_hd__o21a_4
X_1334_ _1330_/Y _1326_/X _1333_/Y VGND VGND VPWR VPWR _1334_/Y sky130_fd_sc_hd__o21ai_4
X_1403_ _1401_/X _1402_/Y VGND VGND VPWR VPWR _2238_/D sky130_fd_sc_hd__nand2_4
XFILLER_51_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1196_ _1193_/X _1194_/X _1195_/Y VGND VGND VPWR VPWR _1196_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_59_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_0_0_m1_clk_local clkbuf_2_1_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_2_0_0_m1_clk_local/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1050_ _1047_/Y _2244_/Q _1048_/X _1049_/Y VGND VGND VPWR VPWR _1060_/A sky130_fd_sc_hd__a22oi_4
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1883_ _1881_/X _1897_/B _2132_/Q VGND VGND VPWR VPWR _1883_/Y sky130_fd_sc_hd__nand3_4
X_1952_ _1952_/A _1083_/A _1952_/C _1952_/D VGND VGND VPWR VPWR _1958_/A sky130_fd_sc_hd__and4_4
XFILLER_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1248_ _1248_/A _1248_/B VGND VGND VPWR VPWR _1248_/Y sky130_fd_sc_hd__nand2_4
X_1317_ _1203_/X _1315_/Y _1344_/B _1366_/B VGND VGND VPWR VPWR _1317_/Y sky130_fd_sc_hd__nand4_4
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1179_ _1176_/Y _1177_/Y _1178_/X VGND VGND VPWR VPWR _1179_/X sky130_fd_sc_hd__o21a_4
XFILLER_24_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2082_ _2073_/CLK _2082_/D VGND VGND VPWR VPWR _2082_/Q sky130_fd_sc_hd__dfxtp_4
X_2220_ _2214_/CLK _1494_/Y VGND VGND VPWR VPWR _1104_/A sky130_fd_sc_hd__dfxtp_4
X_1102_ _2281_/Q _2268_/Q _1101_/X VGND VGND VPWR VPWR _1102_/X sky130_fd_sc_hd__o21a_4
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2151_ _2256_/CLK _1839_/Y VGND VGND VPWR VPWR _2151_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_61_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1033_ _1016_/X VGND VGND VPWR VPWR _1033_/X sky130_fd_sc_hd__buf_2
X_1935_ _1254_/Y _1214_/C _1907_/X _1330_/Y _1934_/X VGND VGND VPWR VPWR _1935_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1797_ _1797_/A VGND VGND VPWR VPWR _1832_/C sky130_fd_sc_hd__buf_2
X_1866_ _1865_/X VGND VGND VPWR VPWR _2140_/D sky130_fd_sc_hd__inv_2
XFILLER_44_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1720_ _1716_/Y _1718_/Y _1719_/X VGND VGND VPWR VPWR _1720_/X sky130_fd_sc_hd__a21o_4
X_1651_ _1651_/A VGND VGND VPWR VPWR _1651_/X sky130_fd_sc_hd__buf_2
X_1582_ _1551_/A _1561_/X _1461_/X VGND VGND VPWR VPWR _1582_/Y sky130_fd_sc_hd__o21ai_4
X_2203_ _2204_/CLK _2203_/D VGND VGND VPWR VPWR _1532_/C sky130_fd_sc_hd__dfxtp_4
X_2065_ _2163_/CLK _1641_/A VGND VGND VPWR VPWR _2059_/D sky130_fd_sc_hd__dfxtp_4
X_2134_ _2133_/CLK _2134_/D VGND VGND VPWR VPWR _1788_/C sky130_fd_sc_hd__dfxtp_4
X_1016_ _1565_/A VGND VGND VPWR VPWR _1016_/X sky130_fd_sc_hd__buf_2
X_1918_ _1757_/A _1879_/D _1918_/C _1918_/D VGND VGND VPWR VPWR _1918_/Y sky130_fd_sc_hd__nand4_4
X_1849_ _1843_/Y _1861_/C _1849_/C VGND VGND VPWR VPWR _1850_/A sky130_fd_sc_hd__and3_4
XFILLER_57_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1634_ _1321_/A VGND VGND VPWR VPWR _1635_/A sky130_fd_sc_hd__buf_2
X_1703_ _1703_/A VGND VGND VPWR VPWR _1704_/B sky130_fd_sc_hd__inv_2
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1565_ _1565_/A VGND VGND VPWR VPWR _1565_/X sky130_fd_sc_hd__buf_2
X_1496_ _1540_/B _1478_/Y _1505_/B _1494_/C VGND VGND VPWR VPWR _2219_/D sky130_fd_sc_hd__and4_4
X_2048_ _2256_/CLK _2053_/Q VGND VGND VPWR VPWR MACRO_RD_SELECT[3] sky130_fd_sc_hd__dfxtp_4
XFILLER_54_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2117_ _2130_/CLK _1917_/Y VGND VGND VPWR VPWR _2015_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1281_ _1192_/Y _1263_/X _1251_/X VGND VGND VPWR VPWR _1281_/X sky130_fd_sc_hd__o21a_4
X_1350_ _1346_/X _1350_/B _1349_/X VGND VGND VPWR VPWR _1350_/Y sky130_fd_sc_hd__nand3_4
XFILLER_48_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1617_ _1617_/A _1560_/B _1613_/A VGND VGND VPWR VPWR _1617_/X sky130_fd_sc_hd__and3_4
X_1548_ _1517_/A _1547_/Y _1542_/X _1539_/A _1074_/X VGND VGND VPWR VPWR _1548_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1479_ _1620_/A _1478_/Y VGND VGND VPWR VPWR _2227_/D sky130_fd_sc_hd__nor2_4
XFILLER_54_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1402_ _1377_/X _2238_/Q VGND VGND VPWR VPWR _1402_/Y sky130_fd_sc_hd__nand2_4
X_1264_ _1264_/A VGND VGND VPWR VPWR _1264_/X sky130_fd_sc_hd__buf_2
X_1333_ _1331_/X _2116_/Q _1410_/A VGND VGND VPWR VPWR _1333_/Y sky130_fd_sc_hd__a21oi_4
X_1195_ _1154_/A _1167_/X _1560_/B VGND VGND VPWR VPWR _1195_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_32_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1882_ _1607_/A VGND VGND VPWR VPWR _1897_/B sky130_fd_sc_hd__buf_2
X_1951_ _1236_/Y _1214_/C _1887_/A _1726_/Y _1934_/X VGND VGND VPWR VPWR _2101_/D
+ sky130_fd_sc_hd__o32ai_4
X_1247_ _1245_/Y _1246_/X VGND VGND VPWR VPWR _1248_/A sky130_fd_sc_hd__nand2_4
X_1178_ _1167_/A VGND VGND VPWR VPWR _1178_/X sky130_fd_sc_hd__buf_2
X_1316_ _1242_/D _1154_/A VGND VGND VPWR VPWR _1344_/B sky130_fd_sc_hd__nor2_4
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1101_ _1101_/A VGND VGND VPWR VPWR _1101_/X sky130_fd_sc_hd__buf_2
X_2150_ _2163_/CLK _1841_/X VGND VGND VPWR VPWR _1838_/B sky130_fd_sc_hd__dfxtp_4
X_1032_ _1028_/Y _1966_/B _1901_/B _1031_/X VGND VGND VPWR VPWR _1032_/X sky130_fd_sc_hd__a211o_4
X_2081_ _2211_/CLK _2089_/Q VGND VGND VPWR VPWR _2081_/Q sky130_fd_sc_hd__dfxtp_4
X_1934_ _1209_/X _1761_/B _1918_/D _1237_/X _1074_/A VGND VGND VPWR VPWR _1934_/X
+ sky130_fd_sc_hd__a41o_4
X_1865_ _1865_/A _1789_/Y VGND VGND VPWR VPWR _1865_/X sky130_fd_sc_hd__xor2_4
X_1796_ _2152_/Q _2151_/Q _1838_/B _1740_/A VGND VGND VPWR VPWR _1797_/A sky130_fd_sc_hd__and4_4
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2279_ _2250_/CLK _2279_/D VGND VGND VPWR VPWR _1030_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_52_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1581_ _1581_/A VGND VGND VPWR VPWR _1581_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1650_ _1237_/X _1835_/A _1918_/D _1318_/X VGND VGND VPWR VPWR _1650_/X sky130_fd_sc_hd__a211o_4
X_2202_ _2027_/CLK _2202_/D VGND VGND VPWR VPWR _2202_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1015_ _1015_/A VGND VGND VPWR VPWR _1565_/A sky130_fd_sc_hd__buf_2
X_2064_ _2028_/CLK _1893_/C VGND VGND VPWR VPWR _2064_/Q sky130_fd_sc_hd__dfxtp_4
X_2133_ _2133_/CLK _1878_/X VGND VGND VPWR VPWR _1876_/B sky130_fd_sc_hd__dfxtp_4
X_1917_ _1236_/Y _1319_/B _1907_/X _1729_/Y _1899_/X VGND VGND VPWR VPWR _1917_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_34_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1779_ _1751_/A _1767_/B _2032_/D VGND VGND VPWR VPWR _1779_/Y sky130_fd_sc_hd__nand3_4
X_1848_ _2148_/Q _1848_/B VGND VGND VPWR VPWR _2148_/D sky130_fd_sc_hd__xnor2_4
XFILLER_8_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_1_0_addressalyzerBlock.SPI_CLK clkbuf_4_1_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2131_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_16_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1564_ _1564_/A _1564_/B _1564_/C _1530_/D VGND VGND VPWR VPWR _1564_/X sky130_fd_sc_hd__and4_4
X_1702_ _2158_/Q _1423_/X _1424_/X _1313_/Y _1318_/X VGND VGND VPWR VPWR _1702_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1633_ _1632_/X _1626_/X _1150_/X _2081_/Q VGND VGND VPWR VPWR _1633_/X sky130_fd_sc_hd__a2bb2o_4
X_1495_ _1494_/B VGND VGND VPWR VPWR _1505_/B sky130_fd_sc_hd__inv_2
XFILLER_62_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2116_ _2124_/CLK _1921_/X VGND VGND VPWR VPWR _2116_/Q sky130_fd_sc_hd__dfxtp_4
X_2047_ _2163_/CLK _2047_/D VGND VGND VPWR VPWR MACRO_RD_SELECT[2] sky130_fd_sc_hd__dfxtp_4
XFILLER_22_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_addressalyzerBlock.SPI_CLK clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1280_ _1279_/Y _1057_/Y _1966_/C _1271_/Y VGND VGND VPWR VPWR _1280_/X sky130_fd_sc_hd__a211o_4
XFILLER_59_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1547_ _1537_/X VGND VGND VPWR VPWR _1547_/Y sky130_fd_sc_hd__inv_2
X_1616_ _1524_/A _1611_/X _2185_/Q VGND VGND VPWR VPWR _1617_/A sky130_fd_sc_hd__a21o_4
X_1478_ _2226_/Q VGND VGND VPWR VPWR _1478_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1401_ _1396_/Y _1397_/Y _1400_/Y VGND VGND VPWR VPWR _1401_/X sky130_fd_sc_hd__a21o_4
X_1263_ _1263_/A VGND VGND VPWR VPWR _1263_/X sky130_fd_sc_hd__buf_2
X_1332_ _1415_/A VGND VGND VPWR VPWR _1410_/A sky130_fd_sc_hd__inv_2
X_1194_ _1156_/A _1156_/B _1185_/Y VGND VGND VPWR VPWR _1194_/X sky130_fd_sc_hd__a21o_4
XFILLER_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1950_ _1301_/Y _1938_/X _1949_/Y VGND VGND VPWR VPWR _2102_/D sky130_fd_sc_hd__o21ai_4
X_1881_ _1897_/A VGND VGND VPWR VPWR _1881_/X sky130_fd_sc_hd__buf_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1315_ _2255_/Q _1152_/A VGND VGND VPWR VPWR _1315_/Y sky130_fd_sc_hd__nor2_4
XFILLER_64_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1246_ _1246_/A VGND VGND VPWR VPWR _1246_/X sky130_fd_sc_hd__buf_2
X_1177_ _2009_/Q _1147_/A VGND VGND VPWR VPWR _1177_/Y sky130_fd_sc_hd__nor2_4
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1100_ _1080_/A _2261_/Q _1099_/X VGND VGND VPWR VPWR _2269_/D sky130_fd_sc_hd__o21a_4
XFILLER_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2080_ _2102_/CLK _2080_/D VGND VGND VPWR VPWR _2080_/Q sky130_fd_sc_hd__dfxtp_4
X_1031_ _2006_/Q _2008_/Q _1029_/A VGND VGND VPWR VPWR _1031_/X sky130_fd_sc_hd__o21a_4
XFILLER_61_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1933_ _1918_/Y _1769_/A _2109_/Q _1349_/X _1932_/Y VGND VGND VPWR VPWR _2109_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_21_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1795_ _1846_/A _1784_/Y _1794_/Y VGND VGND VPWR VPWR _1836_/A sky130_fd_sc_hd__nor3_4
X_1864_ _1864_/A VGND VGND VPWR VPWR _1864_/Y sky130_fd_sc_hd__inv_2
X_2278_ _2250_/CLK _1044_/Y VGND VGND VPWR VPWR _2278_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_37_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1229_ _1229_/A VGND VGND VPWR VPWR _1229_/X sky130_fd_sc_hd__buf_2
XFILLER_57_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1580_ _1564_/B _1564_/A _1579_/Y VGND VGND VPWR VPWR _1581_/A sky130_fd_sc_hd__o21ai_4
XFILLER_7_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2201_ _2204_/CLK _1557_/Y VGND VGND VPWR VPWR _1517_/A sky130_fd_sc_hd__dfxtp_4
X_2132_ _2130_/CLK _1884_/Y VGND VGND VPWR VPWR _2132_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_3_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2063_ _2061_/CLK _2063_/D VGND VGND VPWR VPWR _2063_/Q sky130_fd_sc_hd__dfxtp_4
X_1014_ _1014_/A _1012_/Y _1013_/Y VGND VGND VPWR VPWR _1014_/Y sky130_fd_sc_hd__nand3_4
X_1916_ _1301_/Y _1905_/A _1915_/Y VGND VGND VPWR VPWR _2118_/D sky130_fd_sc_hd__o21ai_4
X_1847_ _1430_/A _1845_/X _1793_/Y _1851_/D VGND VGND VPWR VPWR _1848_/B sky130_fd_sc_hd__nand4_4
X_1778_ _1101_/A _1757_/A _2268_/Q VGND VGND VPWR VPWR _1932_/A sky130_fd_sc_hd__nand3_4
XFILLER_57_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1701_ _1377_/X _1699_/Y _1700_/Y VGND VGND VPWR VPWR _1701_/Y sky130_fd_sc_hd__o21ai_4
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1563_ _2195_/Q VGND VGND VPWR VPWR _1564_/B sky130_fd_sc_hd__buf_2
X_1494_ _1598_/A _1494_/B _1494_/C _1478_/Y VGND VGND VPWR VPWR _1494_/Y sky130_fd_sc_hd__nor4_4
X_1632_ _1344_/Y VGND VGND VPWR VPWR _1632_/X sky130_fd_sc_hd__buf_2
XFILLER_54_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2115_ _2131_/CLK _1925_/Y VGND VGND VPWR VPWR _1411_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_39_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2046_ _2163_/CLK _2051_/Q VGND VGND VPWR VPWR MACRO_RD_SELECT[1] sky130_fd_sc_hd__dfxtp_4
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_5_0_m1_clk_local clkbuf_2_2_0_m1_clk_local/X VGND VGND VPWR VPWR _2187_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1546_ _2204_/Q _1544_/Y _1545_/Y VGND VGND VPWR VPWR _1546_/X sky130_fd_sc_hd__o21a_4
X_1615_ _2186_/Q _1613_/Y _1614_/Y VGND VGND VPWR VPWR _1615_/X sky130_fd_sc_hd__o21a_4
X_1477_ _1620_/A _1080_/X VGND VGND VPWR VPWR _1477_/Y sky130_fd_sc_hd__nor2_4
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2029_ _2256_/CLK _2034_/Q VGND VGND VPWR VPWR MACRO_WR_SELECT[2] sky130_fd_sc_hd__dfxtp_4
XFILLER_10_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1331_ _1325_/A VGND VGND VPWR VPWR _1331_/X sky130_fd_sc_hd__buf_2
X_1400_ _2278_/Q _1398_/X _1630_/B _1400_/D VGND VGND VPWR VPWR _1400_/Y sky130_fd_sc_hd__nand4_4
X_1262_ _1246_/X _1245_/Y _1261_/Y VGND VGND VPWR VPWR _1262_/Y sky130_fd_sc_hd__o21ai_4
X_1193_ _1192_/Y _1177_/Y _1178_/X VGND VGND VPWR VPWR _1193_/X sky130_fd_sc_hd__o21a_4
XFILLER_24_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1529_ _1529_/A VGND VGND VPWR VPWR _1530_/D sky130_fd_sc_hd__inv_2
XFILLER_35_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1880_ _1879_/X VGND VGND VPWR VPWR _1897_/A sky130_fd_sc_hd__inv_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1314_ _1313_/Y VGND VGND VPWR VPWR _1319_/B sky130_fd_sc_hd__buf_2
XFILLER_64_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1176_ _2274_/Q VGND VGND VPWR VPWR _1176_/Y sky130_fd_sc_hd__inv_2
X_1245_ _1245_/A _1057_/Y _1051_/Y _1278_/B VGND VGND VPWR VPWR _1245_/Y sky130_fd_sc_hd__nor4_4
XFILLER_24_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1030_ _1030_/A VGND VGND VPWR VPWR _1901_/B sky130_fd_sc_hd__inv_2
XFILLER_61_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1932_ _1932_/A VGND VGND VPWR VPWR _1932_/Y sky130_fd_sc_hd__inv_2
X_1863_ _1863_/A _1863_/B VGND VGND VPWR VPWR _1864_/A sky130_fd_sc_hd__xor2_4
XFILLER_21_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1794_ _1364_/A _1789_/Y _1857_/D _1793_/Y VGND VGND VPWR VPWR _1794_/Y sky130_fd_sc_hd__nand4_4
X_2277_ _2242_/CLK _2277_/D VGND VGND VPWR VPWR _1071_/B sky130_fd_sc_hd__dfxtp_4
X_1228_ _2249_/Q VGND VGND VPWR VPWR _1229_/A sky130_fd_sc_hd__inv_2
XFILLER_52_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1159_ _1147_/A VGND VGND VPWR VPWR _1217_/A sky130_fd_sc_hd__inv_2
XFILLER_12_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2200_ _2027_/CLK _2200_/D VGND VGND VPWR VPWR _1530_/C sky130_fd_sc_hd__dfxtp_4
X_2131_ _2131_/CLK _2131_/D VGND VGND VPWR VPWR _2131_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_3_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2062_ _2163_/CLK _2126_/Q VGND VGND VPWR VPWR _2056_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_4_6_0_addressalyzerBlock.SPI_CLK clkbuf_4_7_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2268_/CLK sky130_fd_sc_hd__clkbuf_1
X_1013_ _1013_/A VGND VGND VPWR VPWR _1013_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1777_ _1754_/X _1775_/Y _1776_/Y VGND VGND VPWR VPWR _2166_/D sky130_fd_sc_hd__o21ai_4
X_1846_ _1846_/A VGND VGND VPWR VPWR _1851_/D sky130_fd_sc_hd__inv_2
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1915_ _1903_/Y _1940_/B _2118_/Q VGND VGND VPWR VPWR _1915_/Y sky130_fd_sc_hd__nand3_4
XFILLER_25_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1631_ _1627_/Y _1674_/B _1630_/X VGND VGND VPWR VPWR _1631_/Y sky130_fd_sc_hd__o21ai_4
X_1700_ _1722_/A _2175_/Q VGND VGND VPWR VPWR _1700_/Y sky130_fd_sc_hd__nand2_4
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1562_ _1551_/A _1561_/X VGND VGND VPWR VPWR _1564_/A sky130_fd_sc_hd__nor2_4
X_1493_ _1598_/A _1490_/C _1490_/B VGND VGND VPWR VPWR _1493_/Y sky130_fd_sc_hd__nor3_4
XFILLER_39_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2114_ _2124_/CLK _2114_/D VGND VGND VPWR VPWR _2114_/Q sky130_fd_sc_hd__dfxtp_4
X_2045_ _2133_/CLK _2050_/Q VGND VGND VPWR VPWR MACRO_RD_SELECT[0] sky130_fd_sc_hd__dfxtp_4
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1829_ _1319_/A _1829_/B VGND VGND VPWR VPWR _1829_/X sky130_fd_sc_hd__xor2_4
XFILLER_57_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1614_ _1610_/X _1611_/X _2185_/Q _2186_/Q _1565_/X VGND VGND VPWR VPWR _1614_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1545_ _1542_/X _1543_/A _1539_/A _2204_/Q _1074_/X VGND VGND VPWR VPWR _1545_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_5_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1476_ _1476_/A _1473_/Y _1475_/Y VGND VGND VPWR VPWR _2229_/D sky130_fd_sc_hd__nor3_4
XFILLER_35_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2028_ _2028_/CLK _2028_/D VGND VGND VPWR VPWR MACRO_WR_SELECT[1] sky130_fd_sc_hd__dfxtp_4
XFILLER_50_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1330_ _1330_/A VGND VGND VPWR VPWR _1330_/Y sky130_fd_sc_hd__inv_2
X_1261_ _1245_/Y _1246_/X _1966_/C VGND VGND VPWR VPWR _1261_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_51_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1192_ _2272_/Q VGND VGND VPWR VPWR _1192_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1528_ _1528_/A _2198_/Q VGND VGND VPWR VPWR _1529_/A sky130_fd_sc_hd__nand2_4
X_1459_ _1459_/A _1137_/X VGND VGND VPWR VPWR _1459_/X sky130_fd_sc_hd__or2_4
XFILLER_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1244_ _2242_/Q _1244_/B _1054_/A _1244_/D VGND VGND VPWR VPWR _1278_/B sky130_fd_sc_hd__nand4_4
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1313_ _1227_/Y VGND VGND VPWR VPWR _1313_/Y sky130_fd_sc_hd__inv_2
X_1175_ _1168_/Y _1174_/X _1033_/X VGND VGND VPWR VPWR _2255_/D sky130_fd_sc_hd__a21oi_4
XFILLER_32_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1931_ _1301_/Y _1922_/Y _1923_/X _1704_/B _1924_/Y VGND VGND VPWR VPWR _2110_/D
+ sky130_fd_sc_hd__o32ai_4
X_1793_ _1792_/Y VGND VGND VPWR VPWR _1793_/Y sky130_fd_sc_hd__inv_2
X_1862_ _1862_/A _1861_/Y VGND VGND VPWR VPWR _1862_/X sky130_fd_sc_hd__xor2_4
XFILLER_6_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2276_ _2247_/CLK _2276_/D VGND VGND VPWR VPWR _2276_/Q sky130_fd_sc_hd__dfxtp_4
X_1158_ _1645_/A _1152_/Y _1158_/C _1291_/D VGND VGND VPWR VPWR _1158_/Y sky130_fd_sc_hd__nor4_4
X_1227_ _2249_/Q _1918_/C VGND VGND VPWR VPWR _1227_/Y sky130_fd_sc_hd__nor2_4
XFILLER_25_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1089_ _1083_/A VGND VGND VPWR VPWR _1101_/A sky130_fd_sc_hd__buf_2
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_11_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2211_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_7_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2061_ _2061_/CLK _2061_/D VGND VGND VPWR VPWR _2061_/Q sky130_fd_sc_hd__dfxtp_4
X_2130_ _2130_/CLK _2130_/D VGND VGND VPWR VPWR _2066_/D sky130_fd_sc_hd__dfxtp_4
X_1012_ _2005_/Q VGND VGND VPWR VPWR _1012_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1914_ _1294_/Y _1905_/A _1913_/Y VGND VGND VPWR VPWR _2119_/D sky130_fd_sc_hd__o21ai_4
X_1776_ _1767_/A _1767_/B _2166_/Q VGND VGND VPWR VPWR _1776_/Y sky130_fd_sc_hd__nand3_4
X_1845_ _1844_/X VGND VGND VPWR VPWR _1845_/X sky130_fd_sc_hd__buf_2
XFILLER_8_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2259_ _2224_/CLK _1131_/Y VGND VGND VPWR VPWR _2259_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_48_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1630_ _1369_/Y _1630_/B VGND VGND VPWR VPWR _1630_/X sky130_fd_sc_hd__and2_4
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1561_ _1551_/C VGND VGND VPWR VPWR _1561_/X sky130_fd_sc_hd__buf_2
X_1492_ _1492_/A VGND VGND VPWR VPWR _1598_/A sky130_fd_sc_hd__buf_2
X_2044_ _2061_/CLK _2022_/Q VGND VGND VPWR VPWR DATA_TO_HASH[7] sky130_fd_sc_hd__dfxtp_4
X_2113_ _2131_/CLK _2113_/D VGND VGND VPWR VPWR _1638_/A sky130_fd_sc_hd__dfxtp_4
X_1759_ _1754_/X _1607_/X _2171_/Q VGND VGND VPWR VPWR _1759_/Y sky130_fd_sc_hd__nand3_4
X_1828_ _1828_/A _1838_/A _1832_/C _1828_/D VGND VGND VPWR VPWR _1829_/B sky130_fd_sc_hd__nand4_4
XFILLER_45_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1544_ _1543_/Y VGND VGND VPWR VPWR _1544_/Y sky130_fd_sc_hd__inv_2
X_1613_ _1613_/A VGND VGND VPWR VPWR _1613_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1475_ _1138_/X _2229_/Q _1986_/C VGND VGND VPWR VPWR _1475_/Y sky130_fd_sc_hd__a21oi_4
X_2027_ _2027_/CLK _2032_/Q VGND VGND VPWR VPWR MACRO_WR_SELECT[0] sky130_fd_sc_hd__dfxtp_4
XFILLER_35_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1260_ _1253_/X _1258_/Y _1476_/A VGND VGND VPWR VPWR _1260_/Y sky130_fd_sc_hd__a21oi_4
X_1191_ _1187_/X _1190_/Y _1033_/X VGND VGND VPWR VPWR _2253_/D sky130_fd_sc_hd__a21oi_4
XFILLER_36_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_1_0_m1_clk_local clkbuf_2_0_0_m1_clk_local/X VGND VGND VPWR VPWR _2133_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_1527_ _1550_/A _1519_/Y _1520_/Y _1551_/C VGND VGND VPWR VPWR _1530_/B sky130_fd_sc_hd__nor4_4
XFILLER_59_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1389_ _1387_/Y _1336_/X _1388_/Y VGND VGND VPWR VPWR _1389_/Y sky130_fd_sc_hd__o21ai_4
X_1458_ _1456_/Y _1443_/X _1457_/Y VGND VGND VPWR VPWR _1458_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_18_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1243_ _1242_/X VGND VGND VPWR VPWR _1244_/B sky130_fd_sc_hd__buf_2
X_1174_ _1167_/A _1171_/Y _1291_/A VGND VGND VPWR VPWR _1174_/X sky130_fd_sc_hd__a21o_4
X_1312_ _2156_/Q VGND VGND VPWR VPWR _1319_/A sky130_fd_sc_hd__inv_2
XFILLER_2_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1930_ _1294_/Y _1922_/Y _1923_/X _1682_/B _1924_/Y VGND VGND VPWR VPWR _2111_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_14_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1792_ _1673_/C _1857_/A VGND VGND VPWR VPWR _1792_/Y sky130_fd_sc_hd__nand2_4
X_1861_ _1861_/A _1843_/Y _1861_/C _1849_/C VGND VGND VPWR VPWR _1861_/Y sky130_fd_sc_hd__nand4_4
X_2275_ _2075_/CLK _2275_/D VGND VGND VPWR VPWR _2275_/Q sky130_fd_sc_hd__dfxtp_4
X_1157_ _1156_/Y _1242_/D VGND VGND VPWR VPWR _1291_/D sky130_fd_sc_hd__nand2_4
X_1226_ _2248_/Q VGND VGND VPWR VPWR _1918_/C sky130_fd_sc_hd__inv_2
X_1088_ _1080_/X _2266_/Q _1087_/X VGND VGND VPWR VPWR _1088_/X sky130_fd_sc_hd__o21a_4
XFILLER_20_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2060_ _2061_/CLK _2066_/Q VGND VGND VPWR VPWR HASH_ADDR[5] sky130_fd_sc_hd__dfxtp_4
X_1011_ _1005_/A VGND VGND VPWR VPWR _1014_/A sky130_fd_sc_hd__inv_2
XFILLER_19_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1913_ _1903_/Y _1940_/B _1913_/C VGND VGND VPWR VPWR _1913_/Y sky130_fd_sc_hd__nand3_4
X_1775_ _1772_/A _1772_/B _2269_/Q VGND VGND VPWR VPWR _1775_/Y sky130_fd_sc_hd__nand3_4
X_1844_ _1843_/Y _1861_/C _1849_/C _1857_/D VGND VGND VPWR VPWR _1844_/X sky130_fd_sc_hd__and4_4
XFILLER_8_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2258_ _2224_/CLK _1135_/Y VGND VGND VPWR VPWR _1126_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2189_ _2187_/CLK _2189_/D VGND VGND VPWR VPWR _2189_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1209_ _1879_/D VGND VGND VPWR VPWR _1209_/X sky130_fd_sc_hd__buf_2
XFILLER_4_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1560_ _1559_/X _1560_/B _1537_/X VGND VGND VPWR VPWR _2200_/D sky130_fd_sc_hd__and3_4
X_2112_ _2131_/CLK _2112_/D VGND VGND VPWR VPWR _2053_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1491_ _1565_/A VGND VGND VPWR VPWR _1492_/A sky130_fd_sc_hd__buf_2
XFILLER_3_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2043_ _2187_/CLK _2021_/Q VGND VGND VPWR VPWR DATA_TO_HASH[6] sky130_fd_sc_hd__dfxtp_4
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1827_ _1836_/A VGND VGND VPWR VPWR _1838_/A sky130_fd_sc_hd__buf_2
X_1758_ _1115_/X _1772_/B _2274_/Q VGND VGND VPWR VPWR _1758_/Y sky130_fd_sc_hd__nand3_4
X_1689_ _2167_/Q _1689_/B VGND VGND VPWR VPWR _1689_/Y sky130_fd_sc_hd__nand2_4
XFILLER_57_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_2_0_addressalyzerBlock.SPI_CLK clkbuf_2_3_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_5_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1543_ _1543_/A _1542_/X _1539_/A VGND VGND VPWR VPWR _1543_/Y sky130_fd_sc_hd__nand3_4
X_1474_ _1474_/A VGND VGND VPWR VPWR _1986_/C sky130_fd_sc_hd__buf_2
X_1612_ _1610_/X _1611_/X _2185_/Q VGND VGND VPWR VPWR _1613_/A sky130_fd_sc_hd__nand3_4
XFILLER_8_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2026_ _2163_/CLK _2026_/D VGND VGND VPWR VPWR HASH_EN sky130_fd_sc_hd__dfxtp_4
XFILLER_2_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1190_ _1188_/X _1189_/Y _1167_/X VGND VGND VPWR VPWR _1190_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_55_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1526_ _1526_/A _1526_/B _1526_/C _1526_/D VGND VGND VPWR VPWR _1551_/C sky130_fd_sc_hd__nand4_4
X_1457_ _1655_/B _1444_/X _1309_/X VGND VGND VPWR VPWR _1457_/Y sky130_fd_sc_hd__o21ai_4
X_1388_ _1336_/A _2066_/D _1415_/A VGND VGND VPWR VPWR _1388_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_42_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2009_ _2242_/CLK _1985_/Y VGND VGND VPWR VPWR _2009_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_23_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1311_ _1306_/Y _1307_/X _1310_/Y VGND VGND VPWR VPWR _2240_/D sky130_fd_sc_hd__a21oi_4
X_1173_ _1173_/A VGND VGND VPWR VPWR _1291_/A sky130_fd_sc_hd__buf_2
X_1242_ _1156_/Y _1150_/A _1152_/A _1242_/D VGND VGND VPWR VPWR _1242_/X sky130_fd_sc_hd__and4_4
XFILLER_24_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1509_ _2208_/Q VGND VGND VPWR VPWR _1509_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1860_ _1859_/Y VGND VGND VPWR VPWR _1860_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1791_ _1791_/A VGND VGND VPWR VPWR _1857_/D sky130_fd_sc_hd__inv_2
X_2274_ _2075_/CLK _1088_/X VGND VGND VPWR VPWR _2274_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1087_ _1081_/X _2274_/Q _1084_/X VGND VGND VPWR VPWR _1087_/X sky130_fd_sc_hd__o21a_4
XFILLER_52_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1225_ _1986_/D _1147_/X _2269_/Q VGND VGND VPWR VPWR _1225_/Y sky130_fd_sc_hd__o21ai_4
X_1156_ _1156_/A _1156_/B VGND VGND VPWR VPWR _1156_/Y sky130_fd_sc_hd__nor2_4
X_1989_ M1_CLK_IN VGND VGND VPWR VPWR _1989_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1010_ _1005_/A _2005_/Q _1013_/A _1986_/D _1009_/Y VGND VGND VPWR VPWR _1010_/Y
+ sky130_fd_sc_hd__o41ai_4
X_1912_ _1286_/Y _1319_/B _1907_/X _1662_/Y _1899_/X VGND VGND VPWR VPWR _2120_/D
+ sky130_fd_sc_hd__o32ai_4
X_1843_ _1786_/Y _1843_/B _1788_/Y VGND VGND VPWR VPWR _1843_/Y sky130_fd_sc_hd__nor3_4
X_1774_ _1754_/X _1772_/Y _1773_/Y VGND VGND VPWR VPWR _1774_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_57_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2257_ _2224_/CLK _2257_/D VGND VGND VPWR VPWR _1128_/D sky130_fd_sc_hd__dfxtp_4
X_1208_ _1366_/B VGND VGND VPWR VPWR _1879_/D sky130_fd_sc_hd__buf_2
X_2188_ _2027_/CLK _2188_/D VGND VGND VPWR VPWR _1523_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1139_ _1128_/D VGND VGND VPWR VPWR _1139_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1490_ _1540_/B _1490_/B _1490_/C VGND VGND VPWR VPWR _2222_/D sky130_fd_sc_hd__and3_4
XFILLER_3_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2042_ _2027_/CLK _2042_/D VGND VGND VPWR VPWR DATA_TO_HASH[5] sky130_fd_sc_hd__dfxtp_4
X_2111_ _2102_/CLK _2111_/D VGND VGND VPWR VPWR _1681_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_62_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1826_ _1812_/B _1812_/C VGND VGND VPWR VPWR _1826_/X sky130_fd_sc_hd__xor2_4
X_1757_ _1757_/A VGND VGND VPWR VPWR _1772_/B sky130_fd_sc_hd__buf_2
X_1688_ _1326_/X _2095_/Q _1328_/X VGND VGND VPWR VPWR _1688_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1611_ _2184_/Q VGND VGND VPWR VPWR _1611_/X sky130_fd_sc_hd__buf_2
XFILLER_12_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1542_ _2202_/Q VGND VGND VPWR VPWR _1542_/X sky130_fd_sc_hd__buf_2
X_1473_ _1473_/A _1444_/X VGND VGND VPWR VPWR _1473_/Y sky130_fd_sc_hd__nor2_4
XFILLER_54_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2025_ _2256_/CLK _1726_/A VGND VGND VPWR VPWR _2026_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_24_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1809_ _1428_/B _1809_/B _1809_/C _1809_/D VGND VGND VPWR VPWR _1809_/Y sky130_fd_sc_hd__nand4_4
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1387_ _2020_/D VGND VGND VPWR VPWR _1387_/Y sky130_fd_sc_hd__inv_2
X_1525_ _1525_/A _1525_/B _1525_/C _1584_/A VGND VGND VPWR VPWR _1526_/B sky130_fd_sc_hd__nor4_4
X_1456_ _1137_/X _2232_/Q _1455_/X VGND VGND VPWR VPWR _1456_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_19_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2008_ _2211_/CLK _2008_/D VGND VGND VPWR VPWR _2008_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_50_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1310_ _1068_/D _1264_/X _1309_/X VGND VGND VPWR VPWR _1310_/Y sky130_fd_sc_hd__o21ai_4
X_1241_ _1240_/X VGND VGND VPWR VPWR _1241_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1172_ _1150_/A VGND VGND VPWR VPWR _1173_/A sky130_fd_sc_hd__inv_2
XFILLER_17_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1508_ _1508_/A _2210_/Q VGND VGND VPWR VPWR _1508_/Y sky130_fd_sc_hd__nand2_4
XFILLER_46_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1439_ _1439_/A _1439_/B VGND VGND VPWR VPWR _1439_/Y sky130_fd_sc_hd__nand2_4
XFILLER_55_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1790_ _2142_/Q _1861_/A VGND VGND VPWR VPWR _1791_/A sky130_fd_sc_hd__nand2_4
X_2273_ _2075_/CLK _1092_/X VGND VGND VPWR VPWR _2273_/Q sky130_fd_sc_hd__dfxtp_4
X_1224_ _1186_/X _1218_/Y _1219_/X _1220_/Y _1223_/Y VGND VGND VPWR VPWR _2250_/D
+ sky130_fd_sc_hd__a41oi_4
X_1086_ _1080_/X _2267_/Q _1085_/X VGND VGND VPWR VPWR _2275_/D sky130_fd_sc_hd__o21a_4
XFILLER_37_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1155_ _1155_/A _2250_/Q _2249_/Q _2248_/Q VGND VGND VPWR VPWR _1156_/B sky130_fd_sc_hd__nand4_4
X_1988_ EXT_RESET_N_fromHost VGND VGND VPWR VPWR _1988_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_3_0_m1_clk_local clkbuf_2_3_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_2_3_0_m1_clk_local/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_2_0_addressalyzerBlock.SPI_CLK clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR clkbuf_4_5_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_47_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1773_ _1767_/A _1767_/B _2167_/Q VGND VGND VPWR VPWR _1773_/Y sky130_fd_sc_hd__nand3_4
X_1911_ _1192_/Y _1905_/A _1910_/Y VGND VGND VPWR VPWR _2121_/D sky130_fd_sc_hd__o21ai_4
X_1842_ _1740_/X _1838_/A VGND VGND VPWR VPWR _2149_/D sky130_fd_sc_hd__xor2_4
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2256_ _2256_/CLK _1146_/Y VGND VGND VPWR VPWR _2256_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2187_ _2187_/CLK _2187_/D VGND VGND VPWR VPWR _1602_/A sky130_fd_sc_hd__dfxtp_4
X_1207_ _1197_/X VGND VGND VPWR VPWR _1366_/B sky130_fd_sc_hd__inv_2
X_1069_ _1069_/A _1069_/B VGND VGND VPWR VPWR _1069_/Y sky130_fd_sc_hd__nand2_4
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1138_ _1137_/X VGND VGND VPWR VPWR _1138_/X sky130_fd_sc_hd__buf_2
XFILLER_63_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2110_ _2102_/CLK _2110_/D VGND VGND VPWR VPWR _1703_/A sky130_fd_sc_hd__dfxtp_4
X_2041_ _2187_/CLK _2019_/Q VGND VGND VPWR VPWR DATA_TO_HASH[4] sky130_fd_sc_hd__dfxtp_4
XFILLER_62_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1756_ _1751_/X _1920_/A _1755_/Y VGND VGND VPWR VPWR _2172_/D sky130_fd_sc_hd__o21ai_4
X_1825_ _2158_/Q _1825_/B VGND VGND VPWR VPWR _2158_/D sky130_fd_sc_hd__xor2_4
X_1687_ _1683_/X _1686_/X _1339_/X VGND VGND VPWR VPWR _1687_/X sky130_fd_sc_hd__a21o_4
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2239_ _2176_/CLK _2239_/D VGND VGND VPWR VPWR _1378_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_21_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1610_ _1524_/A VGND VGND VPWR VPWR _1610_/X sky130_fd_sc_hd__buf_2
XFILLER_8_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1541_ _1540_/Y VGND VGND VPWR VPWR _2205_/D sky130_fd_sc_hd__inv_2
XFILLER_39_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1472_ _1470_/Y _1972_/A _1471_/Y VGND VGND VPWR VPWR _2230_/D sky130_fd_sc_hd__a21oi_4
XFILLER_54_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2024_ _2101_/CLK _2023_/Q VGND VGND VPWR VPWR _1015_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1739_ _1426_/A _1782_/A _1657_/X VGND VGND VPWR VPWR _1739_/Y sky130_fd_sc_hd__a21oi_4
X_1808_ _1350_/B VGND VGND VPWR VPWR _1810_/A sky130_fd_sc_hd__inv_2
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1524_ _1524_/A _2184_/Q _2185_/Q _2186_/Q VGND VGND VPWR VPWR _1584_/A sky130_fd_sc_hd__nand4_4
X_1386_ _1384_/Y _1336_/X _1385_/Y VGND VGND VPWR VPWR _1386_/Y sky130_fd_sc_hd__o21ai_4
X_1455_ _1127_/X _2233_/Q VGND VGND VPWR VPWR _1455_/X sky130_fd_sc_hd__or2_4
X_2007_ _2247_/CLK _2007_/D VGND VGND VPWR VPWR _1013_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_23_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1240_ _1178_/X _1238_/X _1239_/X VGND VGND VPWR VPWR _1240_/X sky130_fd_sc_hd__a21bo_4
X_1171_ _1152_/Y _1169_/Y _1156_/A _1156_/B _1255_/D VGND VGND VPWR VPWR _1171_/Y
+ sky130_fd_sc_hd__o41ai_4
XFILLER_2_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1507_ _1507_/A VGND VGND VPWR VPWR _1508_/A sky130_fd_sc_hd__inv_2
XFILLER_55_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1438_ _1722_/A _1438_/B VGND VGND VPWR VPWR _1439_/B sky130_fd_sc_hd__nand2_4
X_1369_ _1366_/Y _1227_/Y _1315_/Y _1344_/B _1368_/Y VGND VGND VPWR VPWR _1369_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_11_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2272_ _2075_/CLK _2272_/D VGND VGND VPWR VPWR _2272_/Q sky130_fd_sc_hd__dfxtp_4
X_1223_ _1952_/D _1178_/X _1084_/X VGND VGND VPWR VPWR _1223_/Y sky130_fd_sc_hd__o21ai_4
X_1154_ _1154_/A VGND VGND VPWR VPWR _1156_/A sky130_fd_sc_hd__inv_2
X_1085_ _1081_/X _2275_/Q _1084_/X VGND VGND VPWR VPWR _1085_/X sky130_fd_sc_hd__o21a_4
XFILLER_20_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1987_ _1014_/A _1980_/Y _1986_/Y VGND VGND VPWR VPWR _2008_/D sky130_fd_sc_hd__o21ai_4
XFILLER_20_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1910_ _1903_/Y _1940_/B _1910_/C VGND VGND VPWR VPWR _1910_/Y sky130_fd_sc_hd__nand3_4
XFILLER_19_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1772_ _1772_/A _1772_/B _2270_/Q VGND VGND VPWR VPWR _1772_/Y sky130_fd_sc_hd__nand3_4
X_1841_ _1838_/B _1841_/B VGND VGND VPWR VPWR _1841_/X sky130_fd_sc_hd__xor2_4
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2186_ _2027_/CLK _1615_/X VGND VGND VPWR VPWR _2186_/Q sky130_fd_sc_hd__dfxtp_4
X_2255_ _2242_/CLK _2255_/D VGND VGND VPWR VPWR _2255_/Q sky130_fd_sc_hd__dfxtp_4
X_1206_ _1003_/A _1147_/A _2271_/Q VGND VGND VPWR VPWR _1206_/X sky130_fd_sc_hd__o21a_4
X_1137_ _1137_/A VGND VGND VPWR VPWR _1137_/X sky130_fd_sc_hd__buf_2
X_1068_ _2242_/Q _1067_/X _1068_/C _1068_/D VGND VGND VPWR VPWR _1068_/Y sky130_fd_sc_hd__nand4_4
XFILLER_56_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2040_ _2256_/CLK _2018_/Q VGND VGND VPWR VPWR DATA_TO_HASH[3] sky130_fd_sc_hd__dfxtp_4
XFILLER_47_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1755_ _1754_/X _1607_/X _1755_/C VGND VGND VPWR VPWR _1755_/Y sky130_fd_sc_hd__nand3_4
X_1686_ _1913_/C _1414_/X _1415_/X _1685_/Y VGND VGND VPWR VPWR _1686_/X sky130_fd_sc_hd__a211o_4
XFILLER_30_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1824_ _1816_/D _1816_/B VGND VGND VPWR VPWR _1824_/X sky130_fd_sc_hd__xor2_4
X_2238_ _2176_/CLK _2238_/D VGND VGND VPWR VPWR _2238_/Q sky130_fd_sc_hd__dfxtp_4
X_2169_ _2073_/CLK _1768_/Y VGND VGND VPWR VPWR _2036_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_53_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1540_ _1540_/A _1540_/B _1540_/C VGND VGND VPWR VPWR _1540_/Y sky130_fd_sc_hd__nand3_4
XFILLER_5_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1471_ _1722_/B _1442_/X _1461_/X VGND VGND VPWR VPWR _1471_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_47_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2023_ _2102_/CLK _1988_/Y VGND VGND VPWR VPWR _2023_/Q sky130_fd_sc_hd__dfxtp_4
X_1807_ _1428_/B _1809_/B _1809_/C _1809_/D _1350_/B VGND VGND VPWR VPWR _1807_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1738_ _1645_/A _1736_/Y _1737_/Y VGND VGND VPWR VPWR _1738_/Y sky130_fd_sc_hd__o21ai_4
X_1669_ _1173_/A _2080_/Q _1428_/C _1346_/A VGND VGND VPWR VPWR _1669_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_41_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1523_ _1602_/A _1523_/B VGND VGND VPWR VPWR _1525_/C sky130_fd_sc_hd__nand2_4
X_1454_ _1452_/Y _1443_/X _1453_/Y VGND VGND VPWR VPWR _1454_/Y sky130_fd_sc_hd__a21oi_4
X_1385_ _1331_/X _2114_/Q _1410_/A VGND VGND VPWR VPWR _1385_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_27_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2006_ _2247_/CLK _2006_/D VGND VGND VPWR VPWR _2006_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_51_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1170_ _1213_/A VGND VGND VPWR VPWR _1255_/D sky130_fd_sc_hd__inv_2
XFILLER_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1506_ _2208_/Q _1506_/B VGND VGND VPWR VPWR _1506_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_4_2_0_addressalyzerBlock.SPI_CLK clkbuf_4_3_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2101_/CLK sky130_fd_sc_hd__clkbuf_1
X_1437_ _1432_/Y _1434_/Y _1436_/Y VGND VGND VPWR VPWR _1439_/A sky130_fd_sc_hd__a21o_4
X_1299_ _1295_/B VGND VGND VPWR VPWR _1299_/Y sky130_fd_sc_hd__inv_2
X_1368_ _1360_/Y _1367_/Y VGND VGND VPWR VPWR _1368_/Y sky130_fd_sc_hd__nor2_4
XFILLER_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_7_0_addressalyzerBlock.SPI_CLK clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2271_ _2075_/CLK _1096_/X VGND VGND VPWR VPWR _2271_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_52_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1084_ _1308_/A VGND VGND VPWR VPWR _1084_/X sky130_fd_sc_hd__buf_2
XFILLER_37_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1153_ _1213_/A VGND VGND VPWR VPWR _1158_/C sky130_fd_sc_hd__buf_2
X_1222_ _1936_/B VGND VGND VPWR VPWR _1952_/D sky130_fd_sc_hd__buf_2
XFILLER_52_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1986_ _1607_/X _1986_/B _1986_/C _1986_/D VGND VGND VPWR VPWR _1986_/Y sky130_fd_sc_hd__nand4_4
XFILLER_20_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1840_ _1836_/A _1740_/X VGND VGND VPWR VPWR _1841_/B sky130_fd_sc_hd__and2_4
X_1771_ _1751_/X _1769_/Y _1770_/Y VGND VGND VPWR VPWR _1771_/Y sky130_fd_sc_hd__o21ai_4
X_2254_ _2242_/CLK _1184_/Y VGND VGND VPWR VPWR _1152_/A sky130_fd_sc_hd__dfxtp_4
X_1067_ _1246_/A _2245_/Q _2244_/Q _1048_/X VGND VGND VPWR VPWR _1067_/X sky130_fd_sc_hd__and4_4
X_2185_ _2187_/CLK _1617_/X VGND VGND VPWR VPWR _2185_/Q sky130_fd_sc_hd__dfxtp_4
X_1205_ _1202_/Y _1249_/A _1163_/Y _1249_/C _1360_/C VGND VGND VPWR VPWR _1205_/X
+ sky130_fd_sc_hd__a41o_4
X_1136_ _2219_/Q VGND VGND VPWR VPWR _1137_/A sky130_fd_sc_hd__inv_2
XFILLER_33_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1969_ _1474_/A _1969_/B VGND VGND VPWR VPWR _1969_/Y sky130_fd_sc_hd__nor2_4
XFILLER_56_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1823_ _1822_/Y VGND VGND VPWR VPWR _2160_/D sky130_fd_sc_hd__inv_2
X_1754_ _1751_/A VGND VGND VPWR VPWR _1754_/X sky130_fd_sc_hd__buf_2
X_1685_ _1418_/A _1684_/Y VGND VGND VPWR VPWR _1685_/Y sky130_fd_sc_hd__nor2_4
XFILLER_57_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2237_ _2176_/CLK _1439_/Y VGND VGND VPWR VPWR _1438_/B sky130_fd_sc_hd__dfxtp_4
X_2168_ _2073_/CLK _1771_/Y VGND VGND VPWR VPWR _2035_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_53_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1119_ _2261_/Q _1105_/A _1118_/X VGND VGND VPWR VPWR _1119_/X sky130_fd_sc_hd__o21a_4
X_2099_ _2268_/CLK _1959_/X VGND VGND VPWR VPWR _2099_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1470_ _1137_/X _2229_/Q _1469_/X VGND VGND VPWR VPWR _1470_/Y sky130_fd_sc_hd__o21ai_4
X_2022_ _2061_/CLK _2022_/D VGND VGND VPWR VPWR _2022_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_62_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1806_ _1806_/A VGND VGND VPWR VPWR _1809_/D sky130_fd_sc_hd__inv_2
X_1668_ _1665_/X _1668_/B VGND VGND VPWR VPWR _1668_/Y sky130_fd_sc_hd__nand2_4
X_1599_ _1592_/A _1592_/B _1492_/A VGND VGND VPWR VPWR _1599_/Y sky130_fd_sc_hd__a21oi_4
X_1737_ _1173_/A _2077_/Q _1428_/C _1346_/A VGND VGND VPWR VPWR _1737_/Y sky130_fd_sc_hd__a2bb2oi_4
XFILLER_38_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1522_ _1586_/A VGND VGND VPWR VPWR _1525_/B sky130_fd_sc_hd__inv_2
X_1453_ _2238_/Q _1444_/X _1309_/X VGND VGND VPWR VPWR _1453_/Y sky130_fd_sc_hd__o21ai_4
X_1384_ ID_toHost VGND VGND VPWR VPWR _1384_/Y sky130_fd_sc_hd__inv_2
X_2005_ _2247_/CLK _1971_/X VGND VGND VPWR VPWR _2005_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1505_ _1481_/X _1505_/B VGND VGND VPWR VPWR _1505_/Y sky130_fd_sc_hd__nand2_4
X_1436_ _1398_/X _1747_/A VGND VGND VPWR VPWR _1436_/Y sky130_fd_sc_hd__nand2_4
X_1367_ _1349_/A VGND VGND VPWR VPWR _1367_/Y sky130_fd_sc_hd__inv_2
X_1298_ _1293_/X _1297_/Y _1476_/A VGND VGND VPWR VPWR _1298_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_23_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2270_ _2262_/CLK _2270_/D VGND VGND VPWR VPWR _2270_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_6_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1221_ _1197_/X VGND VGND VPWR VPWR _1936_/B sky130_fd_sc_hd__buf_2
X_1083_ _1083_/A VGND VGND VPWR VPWR _1308_/A sky130_fd_sc_hd__buf_2
X_1152_ _1152_/A VGND VGND VPWR VPWR _1152_/Y sky130_fd_sc_hd__inv_2
X_1985_ _1163_/Y _1984_/Y _1476_/A VGND VGND VPWR VPWR _1985_/Y sky130_fd_sc_hd__a21oi_4
X_1419_ _1905_/C _1414_/X _1415_/X _1418_/Y VGND VGND VPWR VPWR _1419_/X sky130_fd_sc_hd__a211o_4
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1770_ _1767_/A _1767_/B _2035_/D VGND VGND VPWR VPWR _1770_/Y sky130_fd_sc_hd__nand3_4
XFILLER_30_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2184_ _2187_/CLK _1619_/X VGND VGND VPWR VPWR _2184_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2253_ _2250_/CLK _2253_/D VGND VGND VPWR VPWR _1242_/D sky130_fd_sc_hd__dfxtp_4
X_1204_ _1203_/X VGND VGND VPWR VPWR _1360_/C sky130_fd_sc_hd__inv_2
X_1066_ _1046_/Y _1066_/B _1066_/C _1065_/Y VGND VGND VPWR VPWR _1066_/Y sky130_fd_sc_hd__nand4_4
XFILLER_33_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1135_ _1134_/Y VGND VGND VPWR VPWR _1135_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1899_ _1209_/X _1229_/X _1761_/B _1237_/X _1074_/A VGND VGND VPWR VPWR _1899_/X
+ sky130_fd_sc_hd__a41o_4
X_1968_ _2221_/Q VGND VGND VPWR VPWR _1969_/B sky130_fd_sc_hd__inv_2
XFILLER_56_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1753_ _1488_/A _1761_/B _2275_/Q VGND VGND VPWR VPWR _1920_/A sky130_fd_sc_hd__nand3_4
X_1822_ _1809_/C _1809_/B VGND VGND VPWR VPWR _1822_/Y sky130_fd_sc_hd__xnor2_4
X_1684_ _2063_/D VGND VGND VPWR VPWR _1684_/Y sky130_fd_sc_hd__inv_2
X_2167_ _2073_/CLK _1774_/Y VGND VGND VPWR VPWR _2167_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2236_ _2224_/CLK _2236_/D VGND VGND VPWR VPWR _1486_/B sky130_fd_sc_hd__dfxtp_4
X_1118_ _2262_/Q _1104_/A _1115_/X VGND VGND VPWR VPWR _1118_/X sky130_fd_sc_hd__o21a_4
XFILLER_53_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1049_ _2096_/Q VGND VGND VPWR VPWR _1049_/Y sky130_fd_sc_hd__inv_2
X_2098_ _2268_/CLK _2098_/D VGND VGND VPWR VPWR _2098_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_48_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2021_ _2028_/CLK _1905_/C VGND VGND VPWR VPWR _2021_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_50_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1736_ _1732_/Y _1328_/X _1735_/X VGND VGND VPWR VPWR _1736_/Y sky130_fd_sc_hd__a21boi_4
X_1805_ _1394_/B _1805_/B VGND VGND VPWR VPWR _1806_/A sky130_fd_sc_hd__nand2_4
X_1667_ _2035_/D _1689_/B _1328_/X _1666_/Y VGND VGND VPWR VPWR _1668_/B sky130_fd_sc_hd__a211o_4
X_1598_ _1598_/A _1526_/B _1597_/Y VGND VGND VPWR VPWR _1598_/Y sky130_fd_sc_hd__nor3_4
XFILLER_53_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2219_ _2211_/CLK _2219_/D VGND VGND VPWR VPWR _2219_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_14_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1383_ _1326_/X _2098_/Q _1328_/X VGND VGND VPWR VPWR _1383_/Y sky130_fd_sc_hd__a21oi_4
X_1521_ _2189_/Q VGND VGND VPWR VPWR _1525_/A sky130_fd_sc_hd__inv_2
X_1452_ _1125_/X _2234_/Q _1451_/X VGND VGND VPWR VPWR _1452_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_35_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2004_ SCSN_fromHost VGND VGND VPWR VPWR SCSN_toClient sky130_fd_sc_hd__buf_2
XFILLER_23_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_7_0_addressalyzerBlock.SPI_CLK clkbuf_4_7_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2075_/CLK sky130_fd_sc_hd__clkbuf_1
X_1719_ _1788_/C _1361_/Y _1371_/X VGND VGND VPWR VPWR _1719_/X sky130_fd_sc_hd__a21o_4
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1504_ _1481_/X _1490_/B VGND VGND VPWR VPWR _1504_/Y sky130_fd_sc_hd__nand2_4
X_1435_ _2278_/Q VGND VGND VPWR VPWR _1747_/A sky130_fd_sc_hd__buf_2
X_1366_ _1203_/X _1366_/B VGND VGND VPWR VPWR _1366_/Y sky130_fd_sc_hd__nor2_4
XFILLER_62_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1297_ _1296_/Y _1257_/X VGND VGND VPWR VPWR _1297_/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1220_ _1986_/D _1147_/X _2270_/Q VGND VGND VPWR VPWR _1220_/Y sky130_fd_sc_hd__o21ai_4
X_1151_ _1150_/X VGND VGND VPWR VPWR _1645_/A sky130_fd_sc_hd__buf_2
XFILLER_60_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1082_ _1015_/A VGND VGND VPWR VPWR _1083_/A sky130_fd_sc_hd__inv_2
X_1984_ _1986_/C _1147_/X VGND VGND VPWR VPWR _1984_/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1418_ _1418_/A _1418_/B VGND VGND VPWR VPWR _1418_/Y sky130_fd_sc_hd__nor2_4
XFILLER_28_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1349_ _1349_/A VGND VGND VPWR VPWR _1349_/X sky130_fd_sc_hd__buf_2
XFILLER_51_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2183_ _2187_/CLK _1620_/Y VGND VGND VPWR VPWR _1524_/A sky130_fd_sc_hd__dfxtp_4
X_1134_ _1134_/A _1129_/Y _1134_/C VGND VGND VPWR VPWR _1134_/Y sky130_fd_sc_hd__nand3_4
X_2252_ _2250_/CLK _1196_/Y VGND VGND VPWR VPWR _1154_/A sky130_fd_sc_hd__dfxtp_4
X_1203_ _1155_/A VGND VGND VPWR VPWR _1203_/X sky130_fd_sc_hd__buf_2
X_1065_ _1245_/A _2098_/Q _1068_/C _1064_/Y VGND VGND VPWR VPWR _1065_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_33_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1898_ _1932_/A _1881_/X _1897_/Y VGND VGND VPWR VPWR _2125_/D sky130_fd_sc_hd__o21ai_4
X_1967_ _1967_/A _1014_/A _1013_/Y VGND VGND VPWR VPWR _1967_/Y sky130_fd_sc_hd__nand3_4
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1683_ _1947_/C _1414_/X _1410_/X _1682_/Y VGND VGND VPWR VPWR _1683_/X sky130_fd_sc_hd__a211o_4
X_1752_ _1952_/C VGND VGND VPWR VPWR _1761_/B sky130_fd_sc_hd__buf_2
XFILLER_30_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1821_ _1820_/X VGND VGND VPWR VPWR _1821_/Y sky130_fd_sc_hd__inv_2
X_1117_ _2262_/Q _1105_/X _1116_/X VGND VGND VPWR VPWR _2263_/D sky130_fd_sc_hd__o21a_4
X_2166_ _2075_/CLK _2166_/D VGND VGND VPWR VPWR _2166_/Q sky130_fd_sc_hd__dfxtp_4
X_2097_ _2268_/CLK _1961_/X VGND VGND VPWR VPWR _2097_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2235_ _2224_/CLK _2235_/D VGND VGND VPWR VPWR _1447_/B sky130_fd_sc_hd__dfxtp_4
X_1048_ _1048_/A VGND VGND VPWR VPWR _1048_/X sky130_fd_sc_hd__buf_2
XFILLER_21_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2020_ _2027_/CLK _2020_/D VGND VGND VPWR VPWR _2042_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_62_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1666_ _1635_/A _1049_/Y VGND VGND VPWR VPWR _1666_/Y sky130_fd_sc_hd__nor2_4
X_1735_ _2032_/D _1405_/X _1328_/A _1734_/Y VGND VGND VPWR VPWR _1735_/X sky130_fd_sc_hd__a211o_4
XFILLER_7_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1804_ _1819_/A VGND VGND VPWR VPWR _1809_/C sky130_fd_sc_hd__buf_2
X_1597_ _1592_/A _1592_/B _1586_/X VGND VGND VPWR VPWR _1597_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_53_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2149_ _2163_/CLK _2149_/D VGND VGND VPWR VPWR _1740_/A sky130_fd_sc_hd__dfxtp_4
X_2218_ _2211_/CLK _2218_/D VGND VGND VPWR VPWR _1494_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_5_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1520_ _1552_/B VGND VGND VPWR VPWR _1520_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_m1_clk_local clkbuf_0_m1_clk_local/X VGND VGND VPWR VPWR clkbuf_2_3_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_12_0_addressalyzerBlock.SPI_CLK clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2214_/CLK sky130_fd_sc_hd__clkbuf_1
X_1382_ _2170_/Q _1689_/B VGND VGND VPWR VPWR _1382_/Y sky130_fd_sc_hd__nand2_4
X_1451_ _2233_/Q _1137_/X VGND VGND VPWR VPWR _1451_/X sky130_fd_sc_hd__or2_4
XFILLER_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2003_ SCLK_fromHost VGND VGND VPWR VPWR SCLK_toClient sky130_fd_sc_hd__buf_2
XFILLER_50_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1649_ _1798_/B VGND VGND VPWR VPWR _1835_/A sky130_fd_sc_hd__inv_2
X_1718_ _1356_/Y _1862_/A _1361_/Y VGND VGND VPWR VPWR _1718_/Y sky130_fd_sc_hd__a21oi_4
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1503_ _1502_/A MOSI_fromHost VGND VGND VPWR VPWR _1503_/X sky130_fd_sc_hd__and2_4
X_1296_ _1294_/Y _1263_/A _1295_/Y VGND VGND VPWR VPWR _1296_/Y sky130_fd_sc_hd__o21ai_4
X_1365_ _1861_/C VGND VGND VPWR VPWR _1865_/A sky130_fd_sc_hd__inv_2
X_1434_ _1362_/X _1849_/C _1371_/X VGND VGND VPWR VPWR _1434_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_31_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1150_ _1150_/A VGND VGND VPWR VPWR _1150_/X sky130_fd_sc_hd__buf_2
Xclkbuf_3_4_0_m1_clk_local clkbuf_2_2_0_m1_clk_local/X VGND VGND VPWR VPWR _2028_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1081_ _2281_/Q VGND VGND VPWR VPWR _1081_/X sky130_fd_sc_hd__buf_2
X_1983_ _1620_/A _1982_/Y VGND VGND VPWR VPWR _2010_/D sky130_fd_sc_hd__nor2_4
X_1417_ _2131_/Q VGND VGND VPWR VPWR _1418_/B sky130_fd_sc_hd__inv_2
X_1279_ _1279_/A VGND VGND VPWR VPWR _1279_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1348_ _1645_/A _1341_/Y _1347_/Y VGND VGND VPWR VPWR _1348_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_51_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2251_ _2250_/CLK _2251_/D VGND VGND VPWR VPWR _1155_/A sky130_fd_sc_hd__dfxtp_4
X_2182_ _2214_/CLK _2182_/D VGND VGND VPWR VPWR _1069_/B sky130_fd_sc_hd__dfxtp_4
X_1064_ _1064_/A VGND VGND VPWR VPWR _1064_/Y sky130_fd_sc_hd__inv_2
X_1133_ _1125_/X _1126_/B _1128_/D VGND VGND VPWR VPWR _1134_/C sky130_fd_sc_hd__nand3_4
X_1202_ _1201_/X VGND VGND VPWR VPWR _1202_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1966_ _1598_/A _1966_/B _1966_/C VGND VGND VPWR VPWR _2013_/D sky130_fd_sc_hd__nor3_4
X_1897_ _1897_/A _1897_/B _2061_/D VGND VGND VPWR VPWR _1897_/Y sky130_fd_sc_hd__nand3_4
XFILLER_56_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1820_ _1805_/B _1819_/Y VGND VGND VPWR VPWR _1820_/X sky130_fd_sc_hd__xor2_4
X_1751_ _1751_/A VGND VGND VPWR VPWR _1751_/X sky130_fd_sc_hd__buf_2
X_1682_ _1418_/A _1682_/B VGND VGND VPWR VPWR _1682_/Y sky130_fd_sc_hd__nor2_4
XFILLER_38_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2234_ _2224_/CLK _1454_/Y VGND VGND VPWR VPWR _2234_/Q sky130_fd_sc_hd__dfxtp_4
X_2165_ _2075_/CLK _1780_/Y VGND VGND VPWR VPWR _2032_/D sky130_fd_sc_hd__dfxtp_4
X_1116_ _2263_/Q _1106_/X _1115_/X VGND VGND VPWR VPWR _1116_/X sky130_fd_sc_hd__o21a_4
X_1047_ _2097_/Q VGND VGND VPWR VPWR _1047_/Y sky130_fd_sc_hd__inv_2
X_2096_ _2268_/CLK _2096_/D VGND VGND VPWR VPWR _2096_/Q sky130_fd_sc_hd__dfxtp_4
X_1949_ _1945_/A _1954_/B _1949_/C VGND VGND VPWR VPWR _1949_/Y sky130_fd_sc_hd__nand3_4
XFILLER_56_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1803_ _1803_/A _1781_/Y _1812_/B _1812_/C VGND VGND VPWR VPWR _1809_/B sky130_fd_sc_hd__nor4_4
X_1596_ _1587_/X _1526_/B _1595_/Y VGND VGND VPWR VPWR _1596_/X sky130_fd_sc_hd__o21a_4
X_1665_ _1661_/X _1664_/Y _1327_/A VGND VGND VPWR VPWR _1665_/X sky130_fd_sc_hd__a21o_4
X_1734_ _1407_/A _1733_/Y VGND VGND VPWR VPWR _1734_/Y sky130_fd_sc_hd__nor2_4
XFILLER_7_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2217_ _2211_/CLK _2217_/D VGND VGND VPWR VPWR _2217_/Q sky130_fd_sc_hd__dfxtp_4
X_2079_ _2130_/CLK _2087_/Q VGND VGND VPWR VPWR _2079_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2148_ _2133_/CLK _2148_/D VGND VGND VPWR VPWR _2148_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_30_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1450_ _1448_/Y _1443_/X _1449_/Y VGND VGND VPWR VPWR _2235_/D sky130_fd_sc_hd__a21oi_4
X_1381_ _1381_/A _1313_/Y _1318_/X VGND VGND VPWR VPWR _1381_/Y sky130_fd_sc_hd__nor3_4
X_2002_ MOSI_fromHost VGND VGND VPWR VPWR MOSI_toClient sky130_fd_sc_hd__buf_2
XFILLER_35_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1579_ _1564_/A _1564_/B _1492_/A VGND VGND VPWR VPWR _1579_/Y sky130_fd_sc_hd__a21oi_4
X_1717_ _2142_/Q VGND VGND VPWR VPWR _1862_/A sky130_fd_sc_hd__inv_2
X_1648_ _1633_/X _1645_/Y _1647_/Y VGND VGND VPWR VPWR _1648_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_58_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1502_ _1502_/A _2213_/Q VGND VGND VPWR VPWR _2214_/D sky130_fd_sc_hd__and2_4
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1433_ _2139_/Q VGND VGND VPWR VPWR _1849_/C sky130_fd_sc_hd__buf_2
X_1295_ _1058_/Y _1295_/B _1068_/C _1255_/D VGND VGND VPWR VPWR _1295_/Y sky130_fd_sc_hd__nand4_4
X_1364_ _1364_/A VGND VGND VPWR VPWR _1861_/C sky130_fd_sc_hd__buf_2
XFILLER_23_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_addressalyzerBlock.SPI_CLK clkbuf_2_3_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1080_ _1080_/A VGND VGND VPWR VPWR _1080_/X sky130_fd_sc_hd__buf_2
XFILLER_37_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1982_ _2222_/Q _2005_/Q _1972_/A _1147_/X VGND VGND VPWR VPWR _1982_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_9_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1416_ _1324_/A VGND VGND VPWR VPWR _1418_/A sky130_fd_sc_hd__buf_2
X_1347_ _1291_/A _2084_/Q _1428_/C _1346_/X VGND VGND VPWR VPWR _1347_/Y sky130_fd_sc_hd__a2bb2oi_4
XFILLER_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1278_ _1051_/Y _1278_/B VGND VGND VPWR VPWR _1279_/A sky130_fd_sc_hd__nor2_4
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1201_ _1039_/A _1005_/A _1200_/Y VGND VGND VPWR VPWR _1201_/X sky130_fd_sc_hd__o21a_4
X_2250_ _2250_/CLK _2250_/D VGND VGND VPWR VPWR _2250_/Q sky130_fd_sc_hd__dfxtp_4
X_2181_ _2214_/CLK _1622_/X VGND VGND VPWR VPWR _1621_/B sky130_fd_sc_hd__dfxtp_4
X_1063_ _1054_/A VGND VGND VPWR VPWR _1068_/C sky130_fd_sc_hd__buf_2
X_1132_ _1127_/X _1128_/D _1126_/B VGND VGND VPWR VPWR _1134_/A sky130_fd_sc_hd__a21o_4
X_1965_ _1733_/Y _1957_/A _2268_/Q _1958_/A VGND VGND VPWR VPWR _2093_/D sky130_fd_sc_hd__a2bb2o_4
X_1896_ _1651_/X _1775_/Y _1887_/X _1707_/B _1888_/X VGND VGND VPWR VPWR _1896_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_56_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1750_ _1749_/X VGND VGND VPWR VPWR _1751_/A sky130_fd_sc_hd__inv_2
XFILLER_30_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1681_ _1681_/A VGND VGND VPWR VPWR _1682_/B sky130_fd_sc_hd__inv_2
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2233_ _2224_/CLK _1458_/Y VGND VGND VPWR VPWR _2233_/Q sky130_fd_sc_hd__dfxtp_4
X_2164_ _2256_/CLK _2164_/D VGND VGND VPWR VPWR _1350_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_53_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1115_ _1308_/A VGND VGND VPWR VPWR _1115_/X sky130_fd_sc_hd__buf_2
X_2095_ _2268_/CLK _1963_/X VGND VGND VPWR VPWR _2095_/Q sky130_fd_sc_hd__dfxtp_4
X_1046_ _1068_/D _1733_/A VGND VGND VPWR VPWR _1046_/Y sky130_fd_sc_hd__xnor2_4
X_1879_ _1952_/A _1083_/A _1952_/C _1879_/D VGND VGND VPWR VPWR _1879_/X sky130_fd_sc_hd__and4_4
X_1948_ _1294_/Y _1938_/X _1947_/Y VGND VGND VPWR VPWR _2103_/D sky130_fd_sc_hd__o21ai_4
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1733_ _1733_/A VGND VGND VPWR VPWR _1733_/Y sky130_fd_sc_hd__inv_2
X_1802_ _1836_/A _1832_/C _1828_/D _1801_/Y VGND VGND VPWR VPWR _1812_/C sky130_fd_sc_hd__nand4_4
X_1664_ _1662_/Y _1336_/X _1663_/Y VGND VGND VPWR VPWR _1664_/Y sky130_fd_sc_hd__o21ai_4
X_1595_ _1592_/B _1592_/A _1586_/X _1587_/X _1565_/X VGND VGND VPWR VPWR _1595_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_26_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2147_ _2133_/CLK _1852_/X VGND VGND VPWR VPWR _1430_/A sky130_fd_sc_hd__dfxtp_4
X_2216_ _2211_/CLK _1500_/X VGND VGND VPWR VPWR _2216_/Q sky130_fd_sc_hd__dfxtp_4
X_2078_ _2073_/CLK _2078_/D VGND VGND VPWR VPWR _2078_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_14_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1029_ _1029_/A VGND VGND VPWR VPWR _1966_/B sky130_fd_sc_hd__inv_2
XFILLER_30_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1380_ _1798_/A VGND VGND VPWR VPWR _1381_/A sky130_fd_sc_hd__inv_2
X_2001_ EXT_RESET_N_fromHost VGND VGND VPWR VPWR EXT_RESET_N_toClient sky130_fd_sc_hd__buf_2
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1716_ _1702_/Y _1714_/Y _1715_/Y VGND VGND VPWR VPWR _1716_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_58_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1578_ _1520_/Y _1575_/Y _1577_/Y VGND VGND VPWR VPWR _1578_/Y sky130_fd_sc_hd__a21oi_4
X_1647_ _1647_/A _1646_/Y VGND VGND VPWR VPWR _1647_/Y sky130_fd_sc_hd__nor2_4
XFILLER_26_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1363_ _1357_/X _2148_/Q _1362_/X VGND VGND VPWR VPWR _1363_/Y sky130_fd_sc_hd__a21oi_4
X_1432_ _1404_/X _1429_/Y _1431_/Y VGND VGND VPWR VPWR _1432_/Y sky130_fd_sc_hd__o21ai_4
X_1501_ _1502_/A SCLK_fromHost VGND VGND VPWR VPWR _1501_/X sky130_fd_sc_hd__and2_4
X_1294_ _2270_/Q VGND VGND VPWR VPWR _1294_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1981_ _1497_/X _1972_/A _1013_/Y _1967_/A _1980_/Y VGND VGND VPWR VPWR _2006_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_13_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1415_ _1415_/A VGND VGND VPWR VPWR _1415_/X sky130_fd_sc_hd__buf_2
XFILLER_3_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1346_ _1346_/A VGND VGND VPWR VPWR _1346_/X sky130_fd_sc_hd__buf_2
X_1277_ _1273_/Y _1275_/X _1276_/Y VGND VGND VPWR VPWR _1277_/Y sky130_fd_sc_hd__a21oi_4
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2180_ _2124_/CLK _1623_/Y VGND VGND VPWR VPWR _1327_/A sky130_fd_sc_hd__dfxtp_4
X_1200_ _1197_/X _1198_/X _1230_/A VGND VGND VPWR VPWR _1200_/Y sky130_fd_sc_hd__nand3_4
X_1062_ _2245_/Q VGND VGND VPWR VPWR _1245_/A sky130_fd_sc_hd__inv_2
X_1131_ _1124_/Y _1126_/Y _1130_/Y VGND VGND VPWR VPWR _1131_/Y sky130_fd_sc_hd__a21oi_4
X_1895_ _1651_/X _1772_/Y _1887_/X _1684_/Y _1888_/X VGND VGND VPWR VPWR _1895_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1964_ _1064_/Y _1957_/A _2269_/Q _1958_/A VGND VGND VPWR VPWR _1964_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_3_0_0_m1_clk_local clkbuf_2_0_0_m1_clk_local/X VGND VGND VPWR VPWR _2163_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1329_ _1326_/X _1954_/C _1328_/X VGND VGND VPWR VPWR _1329_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1680_ _2103_/Q VGND VGND VPWR VPWR _1947_/C sky130_fd_sc_hd__buf_2
X_1114_ _2263_/Q _1105_/X _1113_/X VGND VGND VPWR VPWR _1114_/X sky130_fd_sc_hd__o21a_4
X_2232_ _2224_/CLK _2232_/D VGND VGND VPWR VPWR _2232_/Q sky130_fd_sc_hd__dfxtp_4
X_2163_ _2163_/CLK _2163_/D VGND VGND VPWR VPWR _1428_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2094_ _2268_/CLK _1964_/X VGND VGND VPWR VPWR _1064_/A sky130_fd_sc_hd__dfxtp_4
X_1045_ _1244_/D VGND VGND VPWR VPWR _1068_/D sky130_fd_sc_hd__buf_2
X_1947_ _1945_/A _1954_/B _1947_/C VGND VGND VPWR VPWR _1947_/Y sky130_fd_sc_hd__nand3_4
X_1878_ _1947_/C _1876_/B VGND VGND VPWR VPWR _1878_/X sky130_fd_sc_hd__xor2_4
XFILLER_56_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1663_ _1331_/X _1893_/C _1415_/X VGND VGND VPWR VPWR _1663_/Y sky130_fd_sc_hd__a21oi_4
X_1732_ _1728_/Y _1732_/B VGND VGND VPWR VPWR _1732_/Y sky130_fd_sc_hd__nand2_4
X_1801_ _1800_/Y VGND VGND VPWR VPWR _1801_/Y sky130_fd_sc_hd__inv_2
X_1594_ _1526_/C _1592_/X _1593_/Y VGND VGND VPWR VPWR _1594_/X sky130_fd_sc_hd__o21a_4
XFILLER_53_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2146_ _2133_/CLK _1855_/X VGND VGND VPWR VPWR _2146_/Q sky130_fd_sc_hd__dfxtp_4
X_2077_ _2176_/CLK _2077_/D VGND VGND VPWR VPWR _2077_/Q sky130_fd_sc_hd__dfxtp_4
X_2215_ _2211_/CLK _1501_/X VGND VGND VPWR VPWR _2215_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1028_ _1028_/A VGND VGND VPWR VPWR _1028_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2000_ VGND VGND VPWR VPWR _2209_/D _2000_/LO sky130_fd_sc_hd__conb_1
XFILLER_35_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_3_0_addressalyzerBlock.SPI_CLK clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR clkbuf_4_7_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_50_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1715_ _1657_/X _1838_/B _1356_/Y VGND VGND VPWR VPWR _1715_/Y sky130_fd_sc_hd__a21oi_4
X_1646_ _1805_/B _1423_/X _1626_/X VGND VGND VPWR VPWR _1646_/Y sky130_fd_sc_hd__nor3_4
X_1577_ _1551_/A _1519_/Y _1520_/Y _1561_/X _1769_/A VGND VGND VPWR VPWR _1577_/Y
+ sky130_fd_sc_hd__o41ai_4
X_2129_ _2131_/CLK _2129_/D VGND VGND VPWR VPWR _1641_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1500_ _1502_/A _2215_/Q VGND VGND VPWR VPWR _1500_/X sky130_fd_sc_hd__and2_4
X_1293_ _1292_/X _1264_/A _1058_/Y VGND VGND VPWR VPWR _1293_/X sky130_fd_sc_hd__a21o_4
X_1431_ _1357_/X _1852_/A _1362_/X VGND VGND VPWR VPWR _1431_/Y sky130_fd_sc_hd__a21oi_4
X_1362_ _1361_/Y VGND VGND VPWR VPWR _1362_/X sky130_fd_sc_hd__buf_2
XFILLER_63_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1629_ _1629_/A VGND VGND VPWR VPWR _1674_/B sky130_fd_sc_hd__buf_2
XFILLER_39_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1980_ _1474_/A _1969_/B _1084_/X VGND VGND VPWR VPWR _1980_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1276_ _2245_/Q _1257_/X _1266_/X VGND VGND VPWR VPWR _1276_/Y sky130_fd_sc_hd__o21ai_4
X_1414_ _1321_/A VGND VGND VPWR VPWR _1414_/X sky130_fd_sc_hd__buf_2
XFILLER_28_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1345_ _1344_/Y VGND VGND VPWR VPWR _1346_/A sky130_fd_sc_hd__inv_2
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1130_ _1999_/C _1129_/Y VGND VGND VPWR VPWR _1130_/Y sky130_fd_sc_hd__nand2_4
X_1061_ _1246_/A _2099_/Q VGND VGND VPWR VPWR _1066_/C sky130_fd_sc_hd__xnor2_4
XFILLER_33_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1894_ _1769_/Y _1881_/X _1893_/Y VGND VGND VPWR VPWR _1894_/Y sky130_fd_sc_hd__o21ai_4
X_1963_ _1055_/Y _1957_/X _2270_/Q _1958_/X VGND VGND VPWR VPWR _1963_/X sky130_fd_sc_hd__a2bb2o_4
X_1328_ _1328_/A VGND VGND VPWR VPWR _1328_/X sky130_fd_sc_hd__buf_2
X_1259_ _1016_/X VGND VGND VPWR VPWR _1476_/A sky130_fd_sc_hd__buf_2
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2231_ _2224_/CLK _2231_/D VGND VGND VPWR VPWR _1459_/A sky130_fd_sc_hd__dfxtp_4
X_1113_ _2264_/Q _1106_/X _1101_/X VGND VGND VPWR VPWR _1113_/X sky130_fd_sc_hd__o21a_4
XFILLER_53_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2093_ _2268_/CLK _2093_/D VGND VGND VPWR VPWR _1733_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_38_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1044_ _1044_/A VGND VGND VPWR VPWR _1044_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2162_ _2256_/CLK _1817_/Y VGND VGND VPWR VPWR _1394_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_46_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1946_ _1286_/Y _1938_/X _1945_/Y VGND VGND VPWR VPWR _1946_/Y sky130_fd_sc_hd__o21ai_4
X_1877_ _1788_/C _1877_/B VGND VGND VPWR VPWR _2134_/D sky130_fd_sc_hd__xnor2_4
XFILLER_29_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1800_ _2156_/Q _1828_/A VGND VGND VPWR VPWR _1800_/Y sky130_fd_sc_hd__nand2_4
X_1662_ _2018_/D VGND VGND VPWR VPWR _1662_/Y sky130_fd_sc_hd__inv_2
X_1731_ _1729_/Y _1331_/X _1730_/Y VGND VGND VPWR VPWR _1732_/B sky130_fd_sc_hd__o21ai_4
XFILLER_7_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2214_ _2214_/CLK _2214_/D VGND VGND VPWR VPWR _2214_/Q sky130_fd_sc_hd__dfxtp_4
X_1593_ _1586_/X _1585_/Y _1587_/X _1526_/C _1565_/X VGND VGND VPWR VPWR _1593_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_53_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2145_ _2133_/CLK _2145_/D VGND VGND VPWR VPWR _1783_/B sky130_fd_sc_hd__dfxtp_4
X_2076_ _2176_/CLK DATA_AVAILABLE[4] VGND VGND VPWR VPWR _2076_/Q sky130_fd_sc_hd__dfxtp_4
X_1027_ _2013_/Q _2011_/Q VGND VGND VPWR VPWR _1028_/A sky130_fd_sc_hd__nor2_4
X_1929_ _1286_/Y _1922_/Y _1923_/X _1659_/Y _1924_/Y VGND VGND VPWR VPWR _2112_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_39_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1576_ _1101_/A VGND VGND VPWR VPWR _1769_/A sky130_fd_sc_hd__buf_2
X_1645_ _1645_/A _1637_/Y _1645_/C VGND VGND VPWR VPWR _1645_/Y sky130_fd_sc_hd__nor3_4
X_1714_ _1709_/X _1712_/Y _1713_/X VGND VGND VPWR VPWR _1714_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_54_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2128_ _2130_/CLK _1894_/Y VGND VGND VPWR VPWR _1893_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_41_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2059_ _2163_/CLK _2059_/D VGND VGND VPWR VPWR HASH_ADDR[4] sky130_fd_sc_hd__dfxtp_4
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1430_ _1430_/A VGND VGND VPWR VPWR _1852_/A sky130_fd_sc_hd__inv_2
XFILLER_36_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1292_ _1295_/B _1068_/C _1158_/C VGND VGND VPWR VPWR _1292_/X sky130_fd_sc_hd__a21o_4
X_1361_ _1200_/Y _1360_/Y VGND VGND VPWR VPWR _1361_/Y sky130_fd_sc_hd__nor2_4
X_1559_ _1552_/A _1564_/C _2199_/Q _1530_/D _1530_/C VGND VGND VPWR VPWR _1559_/X
+ sky130_fd_sc_hd__a41o_4
X_1628_ _1361_/Y VGND VGND VPWR VPWR _1629_/A sky130_fd_sc_hd__inv_2
XFILLER_39_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1413_ _1940_/C _1405_/X _1410_/X _1412_/Y VGND VGND VPWR VPWR _1413_/X sky130_fd_sc_hd__a211o_4
X_1275_ _1274_/Y _1263_/X _1264_/X VGND VGND VPWR VPWR _1275_/X sky130_fd_sc_hd__o21a_4
XFILLER_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1344_ _1315_/Y _1344_/B _1203_/X VGND VGND VPWR VPWR _1344_/Y sky130_fd_sc_hd__nand3_4
XFILLER_59_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1060_ _1060_/A _1060_/B _1056_/Y _1059_/Y VGND VGND VPWR VPWR _1066_/B sky130_fd_sc_hd__and4_4
X_1962_ _1049_/Y _1957_/X _2271_/Q _1958_/X VGND VGND VPWR VPWR _2096_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1893_ _1897_/A _1897_/B _1893_/C VGND VGND VPWR VPWR _1893_/Y sky130_fd_sc_hd__nand3_4
XFILLER_56_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1327_ _1327_/A VGND VGND VPWR VPWR _1328_/A sky130_fd_sc_hd__inv_2
X_1258_ _1258_/A _1257_/X VGND VGND VPWR VPWR _1258_/Y sky130_fd_sc_hd__nand2_4
XFILLER_24_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1189_ _1242_/D _1156_/A _1158_/C _1156_/B VGND VGND VPWR VPWR _1189_/Y sky130_fd_sc_hd__nor4_4
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2230_ _2211_/CLK _2230_/D VGND VGND VPWR VPWR _2230_/Q sky130_fd_sc_hd__dfxtp_4
X_1112_ _2264_/Q _1105_/X _1111_/X VGND VGND VPWR VPWR _1112_/X sky130_fd_sc_hd__o21a_4
XFILLER_38_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2092_ _2131_/CLK DATA_FROM_HASH[7] VGND VGND VPWR VPWR _2084_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1043_ _1038_/X _1041_/Y _1016_/X _1042_/Y VGND VGND VPWR VPWR _1044_/A sky130_fd_sc_hd__a211o_4
X_2161_ _2256_/CLK _1821_/Y VGND VGND VPWR VPWR _1805_/B sky130_fd_sc_hd__dfxtp_4
X_1945_ _1945_/A _1954_/B HASH_LED VGND VGND VPWR VPWR _1945_/Y sky130_fd_sc_hd__nand3_4
XFILLER_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1876_ _1947_/C _1876_/B VGND VGND VPWR VPWR _1877_/B sky130_fd_sc_hd__nand2_4
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_3_0_addressalyzerBlock.SPI_CLK clkbuf_4_3_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2124_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1730_ _1336_/A _2061_/D _1415_/A VGND VGND VPWR VPWR _1730_/Y sky130_fd_sc_hd__a21oi_4
X_1592_ _1592_/A _1592_/B _1586_/X _1587_/X VGND VGND VPWR VPWR _1592_/X sky130_fd_sc_hd__and4_4
X_1661_ HASH_LED _1407_/A _1410_/X _1660_/Y VGND VGND VPWR VPWR _1661_/X sky130_fd_sc_hd__a211o_4
XFILLER_7_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2213_ _2214_/CLK _1503_/X VGND VGND VPWR VPWR _2213_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2144_ _2133_/CLK _1858_/Y VGND VGND VPWR VPWR _1673_/C sky130_fd_sc_hd__dfxtp_4
X_2075_ _2075_/CLK DATA_AVAILABLE[3] VGND VGND VPWR VPWR _2070_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_53_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1026_ _1029_/A _2013_/Q _1026_/C _1026_/D VGND VGND VPWR VPWR _1026_/X sky130_fd_sc_hd__or4_4
X_1928_ _1192_/Y _1922_/Y _1923_/X _1639_/B _1924_/Y VGND VGND VPWR VPWR _2113_/D
+ sky130_fd_sc_hd__o32ai_4
X_1859_ _1857_/A _1845_/X VGND VGND VPWR VPWR _1859_/Y sky130_fd_sc_hd__xnor2_4
Xclkbuf_2_2_0_m1_clk_local clkbuf_2_3_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_2_2_0_m1_clk_local/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1713_ _1423_/X _1424_/X _1150_/A _2078_/Q VGND VGND VPWR VPWR _1713_/X sky130_fd_sc_hd__a2bb2o_4
X_1575_ _1552_/A VGND VGND VPWR VPWR _1575_/Y sky130_fd_sc_hd__inv_2
X_1644_ _1640_/X _1643_/X _1339_/X VGND VGND VPWR VPWR _1645_/C sky130_fd_sc_hd__a21oi_4
X_2127_ _2130_/CLK _1895_/Y VGND VGND VPWR VPWR _2063_/D sky130_fd_sc_hd__dfxtp_4
X_1009_ _1004_/Y _1003_/A _1006_/Y _1008_/Y VGND VGND VPWR VPWR _1009_/Y sky130_fd_sc_hd__a22oi_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2058_ _2028_/CLK _2064_/Q VGND VGND VPWR VPWR HASH_ADDR[3] sky130_fd_sc_hd__dfxtp_4
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1360_ _1315_/Y _1344_/B _1360_/C VGND VGND VPWR VPWR _1360_/Y sky130_fd_sc_hd__nand3_4
X_1291_ _1291_/A _1152_/Y _1290_/Y _1291_/D VGND VGND VPWR VPWR _1295_/B sky130_fd_sc_hd__nor4_4
XFILLER_23_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1558_ _1552_/B VGND VGND VPWR VPWR _1564_/C sky130_fd_sc_hd__buf_2
X_1489_ _1489_/A VGND VGND VPWR VPWR _1490_/B sky130_fd_sc_hd__inv_2
X_1627_ _1627_/A VGND VGND VPWR VPWR _1627_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1412_ _1407_/A _1411_/Y VGND VGND VPWR VPWR _1412_/Y sky130_fd_sc_hd__nor2_4
X_1343_ _1349_/A VGND VGND VPWR VPWR _1428_/C sky130_fd_sc_hd__buf_2
X_1274_ _2273_/Q VGND VGND VPWR VPWR _1274_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1892_ _1651_/X _1765_/Y _1887_/X _1642_/B _1888_/X VGND VGND VPWR VPWR _2129_/D
+ sky130_fd_sc_hd__o32ai_4
X_1961_ _1047_/Y _1957_/X _2272_/Q _1958_/X VGND VGND VPWR VPWR _1961_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_18_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1326_ _1336_/A VGND VGND VPWR VPWR _1326_/X sky130_fd_sc_hd__buf_2
X_1257_ _1264_/A VGND VGND VPWR VPWR _1257_/X sky130_fd_sc_hd__buf_2
X_1188_ _1003_/A _1147_/A _2273_/Q VGND VGND VPWR VPWR _1188_/X sky130_fd_sc_hd__o21a_4
XFILLER_24_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE2_0 EXT_RESET_N_fromHost VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2160_ _2163_/CLK _2160_/D VGND VGND VPWR VPWR _1819_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_61_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1111_ _2265_/Q _1106_/X _1101_/X VGND VGND VPWR VPWR _1111_/X sky130_fd_sc_hd__o21a_4
XFILLER_46_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2091_ _2176_/CLK DATA_FROM_HASH[6] VGND VGND VPWR VPWR _2091_/Q sky130_fd_sc_hd__dfxtp_4
X_1042_ _1035_/X _1038_/B _2278_/Q VGND VGND VPWR VPWR _1042_/Y sky130_fd_sc_hd__a21oi_4
X_1944_ _1192_/Y _1938_/X _1943_/Y VGND VGND VPWR VPWR _2105_/D sky130_fd_sc_hd__o21ai_4
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1875_ _1875_/A VGND VGND VPWR VPWR _1875_/Y sky130_fd_sc_hd__inv_2
X_1309_ _1607_/A VGND VGND VPWR VPWR _1309_/X sky130_fd_sc_hd__buf_2
XFILLER_52_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1660_ _1321_/A _1659_/Y VGND VGND VPWR VPWR _1660_/Y sky130_fd_sc_hd__nor2_4
X_1591_ _2189_/Q VGND VGND VPWR VPWR _1592_/B sky130_fd_sc_hd__buf_2
X_2212_ _2247_/CLK _1504_/Y VGND VGND VPWR VPWR _1490_/C sky130_fd_sc_hd__dfxtp_4
X_2143_ _2133_/CLK _1860_/Y VGND VGND VPWR VPWR _1857_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1025_ _1071_/B _1039_/A _1213_/A _1757_/A VGND VGND VPWR VPWR _1026_/D sky130_fd_sc_hd__a22oi_4
X_2074_ _2102_/CLK DATA_AVAILABLE[2] VGND VGND VPWR VPWR _2074_/Q sky130_fd_sc_hd__dfxtp_4
X_1927_ _1918_/Y _1769_/A _2114_/Q _1349_/X _1926_/Y VGND VGND VPWR VPWR _2114_/D
+ sky130_fd_sc_hd__a32o_4
X_1858_ _1673_/C _1858_/B VGND VGND VPWR VPWR _1858_/Y sky130_fd_sc_hd__xnor2_4
X_1789_ _1785_/Y _1786_/Y _1843_/B _1788_/Y VGND VGND VPWR VPWR _1789_/Y sky130_fd_sc_hd__nor4_4
XFILLER_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1643_ _1910_/C _1635_/A _1415_/X _1642_/Y VGND VGND VPWR VPWR _1643_/X sky130_fd_sc_hd__a211o_4
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1712_ _1710_/Y _1711_/Y _1150_/X VGND VGND VPWR VPWR _1712_/Y sky130_fd_sc_hd__a21oi_4
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1574_ _1528_/A _1530_/B _1573_/Y VGND VGND VPWR VPWR _2197_/D sky130_fd_sc_hd__o21a_4
X_2057_ _2061_/CLK _2063_/Q VGND VGND VPWR VPWR HASH_ADDR[2] sky130_fd_sc_hd__dfxtp_4
X_2126_ _2131_/CLK _1896_/Y VGND VGND VPWR VPWR _2126_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_26_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1008_ _1474_/A _2221_/Q VGND VGND VPWR VPWR _1008_/Y sky130_fd_sc_hd__nor2_4
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1290_ _1244_/D VGND VGND VPWR VPWR _1290_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1626_ _1424_/X VGND VGND VPWR VPWR _1626_/X sky130_fd_sc_hd__buf_2
X_1557_ _1531_/A _1537_/X _1556_/Y VGND VGND VPWR VPWR _1557_/Y sky130_fd_sc_hd__a21oi_4
X_1488_ _1488_/A VGND VGND VPWR VPWR _1540_/B sky130_fd_sc_hd__buf_2
XFILLER_54_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2109_ _2124_/CLK _2109_/D VGND VGND VPWR VPWR _2109_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_27_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1411_ _1411_/A VGND VGND VPWR VPWR _1411_/Y sky130_fd_sc_hd__inv_2
X_1273_ _2245_/Q _1271_/Y _1272_/X VGND VGND VPWR VPWR _1273_/Y sky130_fd_sc_hd__o21ai_4
X_1342_ _1197_/X _1230_/A _1229_/A VGND VGND VPWR VPWR _1349_/A sky130_fd_sc_hd__nor3_4
XFILLER_24_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1609_ _1602_/Y _1584_/X _1608_/Y VGND VGND VPWR VPWR _2187_/D sky130_fd_sc_hd__a21oi_4
XFILLER_59_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1891_ _1761_/Y _1881_/X _1890_/Y VGND VGND VPWR VPWR _2130_/D sky130_fd_sc_hd__o21ai_4
X_1960_ _1052_/Y _1957_/X _2273_/Q _1958_/X VGND VGND VPWR VPWR _2098_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_41_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1325_ _1325_/A VGND VGND VPWR VPWR _1336_/A sky130_fd_sc_hd__buf_2
X_1256_ _1254_/Y _1263_/A _1255_/Y VGND VGND VPWR VPWR _1258_/A sky130_fd_sc_hd__o21ai_4
X_1187_ _1185_/Y _1186_/X _1163_/Y _1249_/C _1169_/Y VGND VGND VPWR VPWR _1187_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_24_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_8_0_addressalyzerBlock.SPI_CLK clkbuf_4_9_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2176_/CLK sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_1 SCLK_fromHost VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2090_ _2073_/CLK DATA_FROM_HASH[5] VGND VGND VPWR VPWR _2082_/D sky130_fd_sc_hd__dfxtp_4
X_1110_ _2265_/Q _1105_/X _1109_/X VGND VGND VPWR VPWR _2266_/D sky130_fd_sc_hd__o21a_4
XFILLER_48_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1041_ _1967_/A _1041_/B _1026_/C VGND VGND VPWR VPWR _1041_/Y sky130_fd_sc_hd__nand3_4
X_1943_ _1945_/A _1940_/B _2105_/Q VGND VGND VPWR VPWR _1943_/Y sky130_fd_sc_hd__nand3_4
X_1874_ _2135_/Q _1873_/Y VGND VGND VPWR VPWR _1875_/A sky130_fd_sc_hd__xor2_4
X_1308_ _1308_/A VGND VGND VPWR VPWR _1607_/A sky130_fd_sc_hd__buf_2
X_1239_ _1237_/X _1167_/A _1101_/A VGND VGND VPWR VPWR _1239_/X sky130_fd_sc_hd__o21a_4
XFILLER_29_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1590_ _1525_/C _1584_/X VGND VGND VPWR VPWR _1592_/A sky130_fd_sc_hd__nor2_4
X_2073_ _2073_/CLK DATA_AVAILABLE[1] VGND VGND VPWR VPWR _2068_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_38_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2211_ _2211_/CLK _1505_/Y VGND VGND VPWR VPWR _1489_/A sky130_fd_sc_hd__dfxtp_4
X_1024_ _1952_/C VGND VGND VPWR VPWR _1757_/A sky130_fd_sc_hd__buf_2
X_2142_ _2133_/CLK _1862_/X VGND VGND VPWR VPWR _2142_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_19_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1926_ _1761_/Y VGND VGND VPWR VPWR _1926_/Y sky130_fd_sc_hd__inv_2
X_1857_ _1857_/A _1789_/Y _1861_/C _1857_/D VGND VGND VPWR VPWR _1858_/B sky130_fd_sc_hd__nand4_4
X_1788_ _2103_/Q _2135_/Q _1788_/C _1876_/B VGND VGND VPWR VPWR _1788_/Y sky130_fd_sc_hd__nand4_4
XFILLER_39_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1642_ _1405_/X _1642_/B VGND VGND VPWR VPWR _1642_/Y sky130_fd_sc_hd__nor2_4
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1711_ _2166_/Q _1689_/B VGND VGND VPWR VPWR _1711_/Y sky130_fd_sc_hd__nand2_4
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1573_ _1564_/B _1564_/A _1564_/C _1528_/A _1565_/X VGND VGND VPWR VPWR _1573_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_3_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2125_ _2073_/CLK _2125_/D VGND VGND VPWR VPWR _2061_/D sky130_fd_sc_hd__dfxtp_4
X_1007_ _1007_/A VGND VGND VPWR VPWR _1474_/A sky130_fd_sc_hd__buf_2
X_2056_ _2163_/CLK _2056_/D VGND VGND VPWR VPWR HASH_ADDR[1] sky130_fd_sc_hd__dfxtp_4
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1909_ _1488_/A VGND VGND VPWR VPWR _1940_/B sky130_fd_sc_hd__buf_2
XFILLER_22_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1556_ _1531_/A _1537_/X _1461_/X VGND VGND VPWR VPWR _1556_/Y sky130_fd_sc_hd__o21ai_4
X_1625_ _1240_/X VGND VGND VPWR VPWR _2178_/D sky130_fd_sc_hd__inv_2
XFILLER_8_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1487_ _1083_/A VGND VGND VPWR VPWR _1488_/A sky130_fd_sc_hd__buf_2
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2108_ _2124_/CLK _1935_/Y VGND VGND VPWR VPWR _1330_/A sky130_fd_sc_hd__dfxtp_4
X_2039_ _2187_/CLK _2017_/Q VGND VGND VPWR VPWR DATA_TO_HASH[2] sky130_fd_sc_hd__dfxtp_4
XFILLER_22_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1410_ _1410_/A VGND VGND VPWR VPWR _1410_/X sky130_fd_sc_hd__buf_2
XFILLER_9_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1272_ _1245_/A _1057_/Y _1051_/Y _1278_/B _1248_/B VGND VGND VPWR VPWR _1272_/X
+ sky130_fd_sc_hd__o41a_4
X_1341_ _1323_/Y _1329_/Y _1340_/Y VGND VGND VPWR VPWR _1341_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_51_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1539_ _1539_/A _1539_/B _2204_/Q CLK_LED VGND VGND VPWR VPWR _1540_/C sky130_fd_sc_hd__nand4_4
X_1608_ _1602_/Y _1584_/X _1607_/X VGND VGND VPWR VPWR _1608_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1890_ _1897_/A _1897_/B _2066_/D VGND VGND VPWR VPWR _1890_/Y sky130_fd_sc_hd__nand3_4
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_13_0_addressalyzerBlock.SPI_CLK clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2262_/CLK sky130_fd_sc_hd__clkbuf_1
X_1255_ _1255_/A _1245_/Y _1246_/X _1255_/D VGND VGND VPWR VPWR _1255_/Y sky130_fd_sc_hd__nand4_4
X_1324_ _1324_/A VGND VGND VPWR VPWR _1325_/A sky130_fd_sc_hd__inv_2
X_1186_ _1249_/A VGND VGND VPWR VPWR _1186_/X sky130_fd_sc_hd__buf_2
XFILLER_64_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XINSDIODE2_2 SCLK_fromHost VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_7_0_m1_clk_local clkbuf_2_3_0_m1_clk_local/X VGND VGND VPWR VPWR _2027_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1040_ _2013_/Q VGND VGND VPWR VPWR _1041_/B sky130_fd_sc_hd__inv_2
X_1942_ _1274_/Y _1214_/C _1907_/X _1384_/Y _1934_/X VGND VGND VPWR VPWR _2106_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1873_ _1947_/C _1788_/C _1876_/B VGND VGND VPWR VPWR _1873_/Y sky130_fd_sc_hd__nand3_4
XFILLER_37_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1307_ _1236_/Y _1263_/A _1251_/X VGND VGND VPWR VPWR _1307_/X sky130_fd_sc_hd__o21a_4
X_1238_ _1236_/Y _1177_/Y _1237_/X _1158_/C VGND VGND VPWR VPWR _1238_/X sky130_fd_sc_hd__o22a_4
X_1169_ _1242_/D VGND VGND VPWR VPWR _1169_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2210_ _2256_/Q _2210_/D SPI_CLK_RESET_N VGND VGND VPWR VPWR _2210_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2072_ _2075_/CLK DATA_AVAILABLE[0] VGND VGND VPWR VPWR _2067_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_53_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2141_ _2133_/CLK _1864_/Y VGND VGND VPWR VPWR _1861_/A sky130_fd_sc_hd__dfxtp_4
X_1023_ _1030_/A VGND VGND VPWR VPWR _1952_/C sky130_fd_sc_hd__buf_2
XFILLER_61_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1925_ _1176_/Y _1922_/Y _1923_/X _1411_/Y _1924_/Y VGND VGND VPWR VPWR _1925_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1787_ _2138_/Q _1627_/A VGND VGND VPWR VPWR _1843_/B sky130_fd_sc_hd__nand2_4
X_1856_ _1854_/A _1794_/Y VGND VGND VPWR VPWR _2145_/D sky130_fd_sc_hd__xor2_4
XFILLER_55_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1572_ _1572_/A VGND VGND VPWR VPWR _1572_/Y sky130_fd_sc_hd__inv_2
X_1641_ _1641_/A VGND VGND VPWR VPWR _1642_/B sky130_fd_sc_hd__inv_2
X_1710_ _1326_/X _1064_/A _1328_/A VGND VGND VPWR VPWR _1710_/Y sky130_fd_sc_hd__a21oi_4
X_2124_ _2124_/CLK _1900_/Y VGND VGND VPWR VPWR _2022_/D sky130_fd_sc_hd__dfxtp_4
X_2055_ _2204_/CLK _2061_/Q VGND VGND VPWR VPWR HASH_ADDR[0] sky130_fd_sc_hd__dfxtp_4
X_1006_ _1006_/A VGND VGND VPWR VPWR _1006_/Y sky130_fd_sc_hd__inv_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1908_ _1274_/Y _1319_/B _1907_/X _1387_/Y _1899_/X VGND VGND VPWR VPWR _1908_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1839_ _2151_/Q _1838_/Y VGND VGND VPWR VPWR _1839_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_1_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1555_ _1554_/Y VGND VGND VPWR VPWR _2202_/D sky130_fd_sc_hd__inv_2
X_1624_ _1186_/X _1218_/Y _1225_/Y _1232_/Y _1234_/Y VGND VGND VPWR VPWR _2179_/D
+ sky130_fd_sc_hd__a41oi_4
XFILLER_54_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2107_ _2131_/CLK _1941_/Y VGND VGND VPWR VPWR _1940_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_39_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1486_ _1502_/A _1486_/B VGND VGND VPWR VPWR _1486_/X sky130_fd_sc_hd__and2_4
XFILLER_54_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2038_ _2163_/CLK _2038_/D VGND VGND VPWR VPWR DATA_TO_HASH[1] sky130_fd_sc_hd__dfxtp_4
X_1340_ _1334_/Y _1338_/Y _1339_/X VGND VGND VPWR VPWR _1340_/Y sky130_fd_sc_hd__a21oi_4
X_1271_ _1271_/A VGND VGND VPWR VPWR _1271_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1538_ _1531_/A _1538_/B _1537_/X VGND VGND VPWR VPWR _1539_/B sky130_fd_sc_hd__nor3_4
X_1607_ _1607_/A VGND VGND VPWR VPWR _1607_/X sky130_fd_sc_hd__buf_2
X_1469_ _2219_/Q _2230_/Q VGND VGND VPWR VPWR _1469_/X sky130_fd_sc_hd__or2_4
XFILLER_50_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1323_ _1755_/C _1689_/B VGND VGND VPWR VPWR _1323_/Y sky130_fd_sc_hd__nand2_4
XFILLER_64_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1254_ _2275_/Q VGND VGND VPWR VPWR _1254_/Y sky130_fd_sc_hd__inv_2
X_1185_ _1156_/A _1156_/B _1255_/D VGND VGND VPWR VPWR _1185_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XINSDIODE2_3 _1913_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1941_ _1176_/Y _1938_/X _1940_/Y VGND VGND VPWR VPWR _1941_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_0_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1872_ _1786_/Y _1788_/Y VGND VGND VPWR VPWR _1872_/X sky130_fd_sc_hd__xor2_4
XFILLER_14_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1306_ _1068_/D _1244_/B _1305_/Y VGND VGND VPWR VPWR _1306_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_64_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1099_ _2281_/Q _2269_/Q _1090_/X VGND VGND VPWR VPWR _1099_/X sky130_fd_sc_hd__o21a_4
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1168_ _1148_/X _1158_/Y _1167_/X VGND VGND VPWR VPWR _1168_/Y sky130_fd_sc_hd__o21ai_4
X_1237_ _1749_/D VGND VGND VPWR VPWR _1237_/X sky130_fd_sc_hd__buf_2
XFILLER_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2140_ _2133_/CLK _2140_/D VGND VGND VPWR VPWR _1364_/A sky130_fd_sc_hd__dfxtp_4
X_2071_ _2176_/CLK _2076_/Q VGND VGND VPWR VPWR _1997_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_19_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1022_ _1022_/A VGND VGND VPWR VPWR _1213_/A sky130_fd_sc_hd__buf_2
XFILLER_61_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1924_ _1918_/Y _1772_/A VGND VGND VPWR VPWR _1924_/Y sky130_fd_sc_hd__nand2_4
X_1855_ _2146_/Q _1854_/Y VGND VGND VPWR VPWR _1855_/X sky130_fd_sc_hd__xor2_4
X_1786_ _1786_/A VGND VGND VPWR VPWR _1786_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2269_ _2262_/CLK _2269_/D VGND VGND VPWR VPWR _2269_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1571_ _1569_/X _1570_/Y VGND VGND VPWR VPWR _1572_/A sky130_fd_sc_hd__nand2_4
X_1640_ _2105_/Q _1635_/A _1410_/X _1639_/Y VGND VGND VPWR VPWR _1640_/X sky130_fd_sc_hd__a211o_4
XFILLER_6_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2123_ _2101_/CLK _1906_/Y VGND VGND VPWR VPWR _1905_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1005_ _1005_/A _1013_/A VGND VGND VPWR VPWR _1006_/A sky130_fd_sc_hd__nor2_4
X_2054_ _2163_/CLK _1638_/A VGND VGND VPWR VPWR _2049_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_19_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1907_ _1887_/A VGND VGND VPWR VPWR _1907_/X sky130_fd_sc_hd__buf_2
X_1838_ _1838_/A _1838_/B _1740_/X VGND VGND VPWR VPWR _1838_/Y sky130_fd_sc_hd__nand3_4
X_1769_ _1769_/A _1772_/B _2271_/Q VGND VGND VPWR VPWR _1769_/Y sky130_fd_sc_hd__nand3_4
XFILLER_1_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1554_ _1542_/X _1543_/A _1553_/Y VGND VGND VPWR VPWR _1554_/Y sky130_fd_sc_hd__o21ai_4
X_1485_ _1485_/A VGND VGND VPWR VPWR _1502_/A sky130_fd_sc_hd__buf_2
X_1623_ _1186_/X _1218_/Y _1219_/X _1220_/Y _1223_/Y VGND VGND VPWR VPWR _1623_/Y
+ sky130_fd_sc_hd__a41oi_4
.ends

