* NGSPICE file created from decred_controller.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

.subckt decred_controller CLK_LED DATA_AVAILABLE DATA_FROM_HASH[0] DATA_FROM_HASH[1]
+ DATA_FROM_HASH[2] DATA_FROM_HASH[3] DATA_FROM_HASH[4] DATA_FROM_HASH[5] DATA_FROM_HASH[6]
+ DATA_FROM_HASH[7] DATA_TO_HASH[0] DATA_TO_HASH[1] DATA_TO_HASH[2] DATA_TO_HASH[3]
+ DATA_TO_HASH[4] DATA_TO_HASH[5] DATA_TO_HASH[6] DATA_TO_HASH[7] EXT_RESET_N_fromHost
+ EXT_RESET_N_toClient HASH_ADDR[0] HASH_ADDR[1] HASH_ADDR[2] HASH_ADDR[3] HASH_ADDR[4]
+ HASH_ADDR[5] HASH_EN HASH_LED ID_fromClient ID_toHost IRQ_OUT_fromClient IRQ_OUT_toHost
+ M1_CLK_IN M1_CLK_SELECT MACRO_RD_SELECT MACRO_WR_SELECT MISO_fromClient MISO_toHost
+ MOSI_fromHost MOSI_toClient PLL_INPUT S1_CLK_IN S1_CLK_SELECT SCLK_fromHost SCLK_toClient
+ SCSN_fromHost SCSN_toClient SPI_CLK_RESET_N THREAD_COUNT[0] THREAD_COUNT[1] THREAD_COUNT[2]
+ THREAD_COUNT[3] m1_clk_local one zero VPWR VGND
XFILLER_54_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2106_ _2108_/CLK _2106_/D VGND VGND VPWR VPWR _1772_/A sky130_fd_sc_hd__dfxtp_4
X_2037_ _2029_/CLK _2037_/D VGND VGND VPWR VPWR _2037_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1270_ _1209_/A VGND VGND VPWR VPWR _1270_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1606_ _1600_/C _1596_/B _1605_/Y VGND VGND VPWR VPWR _2184_/D sky130_fd_sc_hd__o21a_4
XFILLER_59_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1399_ THREAD_COUNT[2] _1421_/A _1397_/Y _1398_/Y VGND VGND VPWR VPWR _1399_/Y sky130_fd_sc_hd__a22oi_4
X_1537_ _2198_/Q _1525_/X _1536_/X VGND VGND VPWR VPWR _2199_/D sky130_fd_sc_hd__o21a_4
X_1468_ _1464_/X _1467_/X _1175_/X VGND VGND VPWR VPWR _1468_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_35_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_m1_clk_local clkbuf_0_m1_clk_local/X VGND VGND VPWR VPWR clkbuf_2_1_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
X_1322_ _1322_/A VGND VGND VPWR VPWR _1323_/C sky130_fd_sc_hd__buf_2
X_1253_ _1253_/A _1155_/X VGND VGND VPWR VPWR _1253_/Y sky130_fd_sc_hd__nand2_4
XFILLER_64_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1184_ _1184_/A _1048_/D _1218_/A VGND VGND VPWR VPWR _1185_/A sky130_fd_sc_hd__nor3_4
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1940_ _1765_/Y VGND VGND VPWR VPWR _1940_/Y sky130_fd_sc_hd__inv_2
X_1871_ _1864_/Y VGND VGND VPWR VPWR _1871_/X sky130_fd_sc_hd__buf_2
XFILLER_9_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_0_m1_clk_local m1_clk_local VGND VGND VPWR VPWR clkbuf_0_m1_clk_local/X sky130_fd_sc_hd__clkbuf_16
X_1236_ _1236_/A VGND VGND VPWR VPWR _1236_/Y sky130_fd_sc_hd__inv_2
X_1305_ _1917_/A VGND VGND VPWR VPWR _1675_/B sky130_fd_sc_hd__buf_2
XFILLER_52_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1098_ _1098_/A VGND VGND VPWR VPWR _1098_/X sky130_fd_sc_hd__buf_2
X_1167_ _1164_/X _2076_/Q _1166_/X VGND VGND VPWR VPWR _1167_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_20_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_m1_clk_local clkbuf_3_3_0_m1_clk_local/A VGND VGND VPWR VPWR _2124_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_2070_ _2213_/CLK _2070_/D VGND VGND VPWR VPWR _2070_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1021_ _1024_/A _0996_/X _1020_/X VGND VGND VPWR VPWR _1021_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_19_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1785_ _2124_/Q _1813_/A VGND VGND VPWR VPWR _1785_/Y sky130_fd_sc_hd__nand2_4
X_1854_ _1371_/X _1774_/D VGND VGND VPWR VPWR _1854_/Y sky130_fd_sc_hd__nor2_4
X_1923_ _1902_/Y _1916_/X _1922_/Y VGND VGND VPWR VPWR _1923_/Y sky130_fd_sc_hd__o21ai_4
X_1219_ _1201_/B _1219_/B VGND VGND VPWR VPWR _1344_/A sky130_fd_sc_hd__nor2_4
X_2199_ _2194_/CLK _2199_/D VGND VGND VPWR VPWR _2199_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1570_ _1570_/A SPI_CLK_RESET_N _1570_/C _1569_/X VGND VGND VPWR VPWR _2189_/D sky130_fd_sc_hd__and4_4
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2122_ _2025_/CLK _1818_/Y VGND VGND VPWR VPWR _2122_/Q sky130_fd_sc_hd__dfxtp_4
X_2053_ _2044_/CLK DATA_FROM_HASH[0] VGND VGND VPWR VPWR _2053_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1004_ _1004_/A VGND VGND VPWR VPWR _1004_/X sky130_fd_sc_hd__buf_2
XFILLER_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1837_ _2115_/Q _1836_/Y VGND VGND VPWR VPWR _1837_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_30_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1768_ _1746_/A _1765_/Y _1767_/Y VGND VGND VPWR VPWR _2133_/D sky130_fd_sc_hd__o21ai_4
X_1906_ _1904_/Y _1473_/B _1905_/X _1407_/Y _1889_/X VGND VGND VPWR VPWR _2086_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_57_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1699_ _1697_/A _2149_/Q VGND VGND VPWR VPWR _1699_/X sky130_fd_sc_hd__and2_4
XFILLER_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1622_ _1621_/C _1608_/Y _1587_/A _1587_/D _1102_/A VGND VGND VPWR VPWR _1622_/Y
+ sky130_fd_sc_hd__a41oi_4
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1484_ _1059_/B _1484_/B VGND VGND VPWR VPWR _1484_/X sky130_fd_sc_hd__xor2_4
X_1553_ _2158_/Q VGND VGND VPWR VPWR _1553_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2105_ _2115_/CLK _1855_/X VGND VGND VPWR VPWR _2105_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2036_ _2171_/CLK _2036_/D VGND VGND VPWR VPWR HASH_ADDR[5] sky130_fd_sc_hd__dfxtp_4
XFILLER_62_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1605_ _1574_/A _1604_/Y _1600_/B _1600_/C _1102_/A VGND VGND VPWR VPWR _1605_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1536_ _2199_/Q _1526_/X _1535_/X VGND VGND VPWR VPWR _1536_/X sky130_fd_sc_hd__o21a_4
X_1398_ _1773_/B _1397_/B _1344_/A _1708_/A VGND VGND VPWR VPWR _1398_/Y sky130_fd_sc_hd__a2bb2oi_4
XFILLER_27_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1467_ _2001_/D _1355_/X _1172_/X _1466_/Y VGND VGND VPWR VPWR _1467_/X sky130_fd_sc_hd__a211o_4
X_2019_ _2171_/CLK _2019_/D VGND VGND VPWR VPWR MACRO_WR_SELECT sky130_fd_sc_hd__dfxtp_4
XFILLER_6_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1252_ _1252_/A _1251_/Y VGND VGND VPWR VPWR _2231_/D sky130_fd_sc_hd__nand2_4
X_1321_ _1971_/A _1971_/B _1064_/Y _1066_/D _1001_/A VGND VGND VPWR VPWR _1322_/A
+ sky130_fd_sc_hd__a41o_4
XFILLER_64_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1183_ _1047_/A VGND VGND VPWR VPWR _1218_/A sky130_fd_sc_hd__inv_2
XFILLER_17_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_4_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_4_9_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
X_1519_ _2215_/Q _1133_/X _1510_/X VGND VGND VPWR VPWR _1519_/X sky130_fd_sc_hd__o21a_4
XFILLER_55_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1870_ _1930_/A _1865_/X _1869_/Y VGND VGND VPWR VPWR _2099_/D sky130_fd_sc_hd__o21ai_4
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1304_ _1005_/Y VGND VGND VPWR VPWR _1917_/A sky130_fd_sc_hd__buf_2
X_1166_ _1166_/A VGND VGND VPWR VPWR _1166_/X sky130_fd_sc_hd__buf_2
X_1235_ _1232_/Y _1233_/X _1234_/Y VGND VGND VPWR VPWR _1235_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_64_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1097_ _1097_/A VGND VGND VPWR VPWR _1097_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1999_ _2182_/CLK _1383_/A VGND VGND VPWR VPWR _1999_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1020_ _1020_/A _1020_/B VGND VGND VPWR VPWR _1020_/X sky130_fd_sc_hd__or2_4
XFILLER_19_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1922_ _1915_/Y _1917_/X _1857_/A VGND VGND VPWR VPWR _1922_/Y sky130_fd_sc_hd__nand3_4
X_1784_ _1783_/Y VGND VGND VPWR VPWR _1815_/C sky130_fd_sc_hd__inv_2
X_1853_ _1772_/A _1853_/B VGND VGND VPWR VPWR _2106_/D sky130_fd_sc_hd__xor2_4
XFILLER_6_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1149_ _1149_/A _1149_/B VGND VGND VPWR VPWR _1182_/B sky130_fd_sc_hd__nor2_4
XFILLER_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1218_ _1218_/A VGND VGND VPWR VPWR _1219_/B sky130_fd_sc_hd__buf_2
X_2198_ _2194_/CLK _2198_/D VGND VGND VPWR VPWR _2198_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_52_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2052_ _2052_/CLK _2052_/D VGND VGND VPWR VPWR _1180_/A sky130_fd_sc_hd__dfxtp_4
X_2121_ _2025_/CLK _1820_/X VGND VGND VPWR VPWR _2121_/Q sky130_fd_sc_hd__dfxtp_4
X_1003_ _1003_/A VGND VGND VPWR VPWR _1003_/X sky130_fd_sc_hd__buf_2
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1905_ _1887_/Y VGND VGND VPWR VPWR _1905_/X sky130_fd_sc_hd__buf_2
X_1836_ _1847_/B _1776_/Y _1832_/C _1832_/D VGND VGND VPWR VPWR _1836_/Y sky130_fd_sc_hd__nand4_4
XFILLER_30_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1767_ _1738_/Y _1767_/B _1767_/C VGND VGND VPWR VPWR _1767_/Y sky130_fd_sc_hd__nand3_4
X_1698_ _1697_/A SCLK_fromHost VGND VGND VPWR VPWR _1698_/X sky130_fd_sc_hd__and2_4
XFILLER_57_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1621_ _1619_/Y _1621_/B _1621_/C _1587_/D VGND VGND VPWR VPWR _1621_/X sky130_fd_sc_hd__and4_4
X_1552_ _1551_/X VGND VGND VPWR VPWR _2194_/D sky130_fd_sc_hd__inv_2
X_2104_ _2115_/CLK _1856_/X VGND VGND VPWR VPWR _1370_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_39_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1483_ _1105_/B _1483_/B VGND VGND VPWR VPWR _1483_/X sky130_fd_sc_hd__xor2_4
X_2035_ _2025_/CLK _2041_/Q VGND VGND VPWR VPWR HASH_ADDR[4] sky130_fd_sc_hd__dfxtp_4
X_1819_ _1827_/B _1815_/B VGND VGND VPWR VPWR _1819_/Y sky130_fd_sc_hd__nand2_4
XFILLER_45_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1604_ _1604_/A VGND VGND VPWR VPWR _1604_/Y sky130_fd_sc_hd__inv_2
X_1535_ _1625_/A VGND VGND VPWR VPWR _1535_/X sky130_fd_sc_hd__buf_2
X_1397_ _1397_/A _1397_/B _1397_/C VGND VGND VPWR VPWR _1397_/Y sky130_fd_sc_hd__nand3_4
X_1466_ _1412_/A _1466_/B VGND VGND VPWR VPWR _1466_/Y sky130_fd_sc_hd__nor2_4
X_2018_ _2124_/CLK _2017_/Q VGND VGND VPWR VPWR HASH_EN sky130_fd_sc_hd__dfxtp_4
XFILLER_42_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1320_ _1449_/B VGND VGND VPWR VPWR _1971_/B sky130_fd_sc_hd__inv_2
XFILLER_64_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1251_ _1274_/A _2231_/Q VGND VGND VPWR VPWR _1251_/Y sky130_fd_sc_hd__nand2_4
X_1182_ _1148_/A _1182_/B _1182_/C VGND VGND VPWR VPWR _1189_/A sky130_fd_sc_hd__nand3_4
XFILLER_64_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1449_ _2010_/Q _1449_/B _1449_/C VGND VGND VPWR VPWR _1449_/Y sky130_fd_sc_hd__nor3_4
X_1518_ _1501_/Y _2198_/Q _1517_/X VGND VGND VPWR VPWR _1518_/X sky130_fd_sc_hd__o21a_4
XFILLER_23_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1303_ _1112_/A _1279_/Y _1291_/A _1302_/Y VGND VGND VPWR VPWR _1307_/A sky130_fd_sc_hd__a211o_4
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1096_ _1894_/A _1078_/X _1079_/X VGND VGND VPWR VPWR _1096_/Y sky130_fd_sc_hd__a21oi_4
X_1234_ _1164_/X _2075_/Q _1166_/A VGND VGND VPWR VPWR _1234_/Y sky130_fd_sc_hd__a21oi_4
X_1165_ _2143_/Q VGND VGND VPWR VPWR _1166_/A sky130_fd_sc_hd__inv_2
XFILLER_20_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1998_ _2189_/CLK _1998_/D VGND VGND VPWR VPWR _1998_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_18_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1852_ _1477_/Y _1371_/X _1774_/D VGND VGND VPWR VPWR _1853_/B sky130_fd_sc_hd__nor3_4
X_1921_ _1316_/Y _1916_/X _1920_/Y VGND VGND VPWR VPWR _2080_/D sky130_fd_sc_hd__o21ai_4
X_1783_ _2122_/Q _2121_/Q VGND VGND VPWR VPWR _1783_/Y sky130_fd_sc_hd__nand2_4
XFILLER_57_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1217_ _1217_/A VGND VGND VPWR VPWR _1217_/X sky130_fd_sc_hd__buf_2
X_1148_ _1148_/A VGND VGND VPWR VPWR _1344_/C sky130_fd_sc_hd__buf_2
X_1079_ _1067_/Y VGND VGND VPWR VPWR _1079_/X sky130_fd_sc_hd__buf_2
XFILLER_25_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2197_ _2194_/CLK _1541_/X VGND VGND VPWR VPWR _2197_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_4_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2120_ _2025_/CLK _1822_/X VGND VGND VPWR VPWR _2120_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2051_ _2051_/CLK _2059_/Q VGND VGND VPWR VPWR _1241_/A sky130_fd_sc_hd__dfxtp_4
X_1002_ _1004_/A VGND VGND VPWR VPWR _1003_/A sky130_fd_sc_hd__buf_2
XFILLER_34_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1835_ _1835_/A VGND VGND VPWR VPWR _1847_/B sky130_fd_sc_hd__buf_2
X_1904_ _1904_/A VGND VGND VPWR VPWR _1904_/Y sky130_fd_sc_hd__inv_2
X_1766_ _1008_/A VGND VGND VPWR VPWR _1767_/B sky130_fd_sc_hd__buf_2
X_1697_ _1697_/A _2151_/Q VGND VGND VPWR VPWR _2152_/D sky130_fd_sc_hd__and2_4
XFILLER_40_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1620_ _1576_/A VGND VGND VPWR VPWR _1621_/B sky130_fd_sc_hd__buf_2
X_1482_ _1482_/A _1126_/B VGND VGND VPWR VPWR _1482_/Y sky130_fd_sc_hd__nor2_4
XFILLER_8_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1551_ _1455_/C _1549_/Y _1550_/Y VGND VGND VPWR VPWR _1551_/X sky130_fd_sc_hd__a21o_4
X_2103_ _2108_/CLK _2103_/D VGND VGND VPWR VPWR _1773_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_39_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2034_ _2029_/CLK _2034_/D VGND VGND VPWR VPWR HASH_ADDR[3] sky130_fd_sc_hd__dfxtp_4
XFILLER_22_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1818_ _2122_/Q _1817_/Y VGND VGND VPWR VPWR _1818_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1749_ _1738_/Y VGND VGND VPWR VPWR _1754_/A sky130_fd_sc_hd__buf_2
XFILLER_45_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_4_0_addressalyzerBlock.SPI_CLK clkbuf_4_5_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2051_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_13_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1603_ _2185_/Q _1601_/Y _1602_/Y VGND VGND VPWR VPWR _2185_/D sky130_fd_sc_hd__o21a_4
XFILLER_4_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1534_ _2199_/Q _1525_/X _1533_/X VGND VGND VPWR VPWR _2200_/D sky130_fd_sc_hd__o21a_4
X_1465_ _2041_/D VGND VGND VPWR VPWR _1466_/B sky130_fd_sc_hd__inv_2
X_2017_ _2124_/CLK _2017_/D VGND VGND VPWR VPWR _2017_/Q sky130_fd_sc_hd__dfxtp_4
X_1396_ _1396_/A _1843_/A _1396_/C VGND VGND VPWR VPWR _1397_/C sky130_fd_sc_hd__nand3_4
XFILLER_12_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1250_ _1246_/Y _1247_/Y _1249_/X VGND VGND VPWR VPWR _1252_/A sky130_fd_sc_hd__a21o_4
XFILLER_49_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1181_ _1088_/X _1177_/Y _1180_/X VGND VGND VPWR VPWR _1181_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_32_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1448_ _1448_/A _1451_/B _1451_/C VGND VGND VPWR VPWR _1448_/Y sky130_fd_sc_hd__nor3_4
X_1517_ _2215_/Q _1902_/A _1510_/X VGND VGND VPWR VPWR _1517_/X sky130_fd_sc_hd__o21a_4
X_1379_ _1773_/A VGND VGND VPWR VPWR _1857_/A sky130_fd_sc_hd__buf_2
XFILLER_46_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1302_ _1086_/X _1049_/X _1296_/Y VGND VGND VPWR VPWR _1302_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1233_ _1170_/A VGND VGND VPWR VPWR _1233_/X sky130_fd_sc_hd__buf_2
XFILLER_64_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1095_ _1748_/C VGND VGND VPWR VPWR _1894_/A sky130_fd_sc_hd__buf_2
X_1164_ _1170_/A VGND VGND VPWR VPWR _1164_/X sky130_fd_sc_hd__buf_2
XFILLER_60_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1997_ _2108_/CLK _1997_/D VGND VGND VPWR VPWR _1997_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_20_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_addressalyzerBlock.SPI_CLK clkbuf_0_addressalyzerBlock.SPI_CLK/X VGND
+ VGND VPWR VPWR clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_7_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1851_ _1834_/C _1834_/A VGND VGND VPWR VPWR _1851_/X sky130_fd_sc_hd__xor2_4
X_1920_ _1915_/Y _1917_/X HASH_LED VGND VGND VPWR VPWR _1920_/Y sky130_fd_sc_hd__nand3_4
X_1782_ _1782_/A VGND VGND VPWR VPWR _1815_/B sky130_fd_sc_hd__buf_2
XFILLER_6_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1216_ _1226_/A _1215_/Y VGND VGND VPWR VPWR _1223_/A sky130_fd_sc_hd__nor2_4
X_2196_ _2194_/CLK _1543_/X VGND VGND VPWR VPWR _2196_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_52_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1147_ _1178_/A _1147_/B VGND VGND VPWR VPWR _1148_/A sky130_fd_sc_hd__nor2_4
X_1078_ _2012_/Q VGND VGND VPWR VPWR _1078_/X sky130_fd_sc_hd__buf_2
XFILLER_25_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2050_ _2058_/CLK _2050_/D VGND VGND VPWR VPWR _1263_/A sky130_fd_sc_hd__dfxtp_4
X_1001_ _1001_/A VGND VGND VPWR VPWR _1004_/A sky130_fd_sc_hd__inv_2
XFILLER_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1834_ _1834_/A _1834_/B _1834_/C VGND VGND VPWR VPWR _1835_/A sky130_fd_sc_hd__and3_4
X_1765_ _1633_/A _1740_/X _2204_/Q VGND VGND VPWR VPWR _1765_/Y sky130_fd_sc_hd__nand3_4
X_1903_ _1902_/Y _1885_/X _1888_/X _1383_/Y _1890_/X VGND VGND VPWR VPWR _2087_/D
+ sky130_fd_sc_hd__o32ai_4
X_1696_ _1694_/X SCSN_fromHost VGND VGND VPWR VPWR _1696_/X sky130_fd_sc_hd__or2_4
X_2248_ _2248_/CLK _1990_/Y VGND VGND VPWR VPWR _1987_/A sky130_fd_sc_hd__dfxtp_4
X_2179_ _2182_/CLK _2179_/D VGND VGND VPWR VPWR _1627_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_40_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1481_ _1479_/X _1223_/A _1480_/X VGND VGND VPWR VPWR _1481_/X sky130_fd_sc_hd__a21o_4
X_1550_ _1455_/C _1549_/Y _1456_/Y VGND VGND VPWR VPWR _1550_/Y sky130_fd_sc_hd__o21ai_4
X_2102_ _2108_/CLK _1861_/Y VGND VGND VPWR VPWR _2102_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2033_ _2182_/CLK _2033_/D VGND VGND VPWR VPWR HASH_ADDR[2] sky130_fd_sc_hd__dfxtp_4
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1817_ _1827_/B _2121_/Q _1815_/B VGND VGND VPWR VPWR _1817_/Y sky130_fd_sc_hd__nand3_4
XFILLER_30_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1748_ _1633_/A _1740_/X _1748_/C VGND VGND VPWR VPWR _1748_/Y sky130_fd_sc_hd__nand3_4
X_1679_ _1679_/A VGND VGND VPWR VPWR _1693_/B sky130_fd_sc_hd__inv_2
XFILLER_38_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1602_ _1600_/B _1589_/B _1600_/C _2185_/Q _1102_/A VGND VGND VPWR VPWR _1602_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_8_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1395_ _1378_/Y _1393_/Y _1394_/X VGND VGND VPWR VPWR _1397_/A sky130_fd_sc_hd__o21ai_4
X_1533_ _2200_/Q _1526_/X _1521_/X VGND VGND VPWR VPWR _1533_/X sky130_fd_sc_hd__o21a_4
X_1464_ _2081_/Q _1355_/X _1166_/X _1463_/Y VGND VGND VPWR VPWR _1464_/X sky130_fd_sc_hd__a211o_4
X_2016_ _2248_/CLK _1975_/X VGND VGND VPWR VPWR _1448_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_50_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1180_ _1180_/A _1179_/X VGND VGND VPWR VPWR _1180_/X sky130_fd_sc_hd__or2_4
XFILLER_17_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1516_ _1501_/Y _2199_/Q _1515_/X VGND VGND VPWR VPWR _1516_/X sky130_fd_sc_hd__o21a_4
X_1378_ _1788_/A _1243_/B _1243_/C _1473_/B _1473_/C VGND VGND VPWR VPWR _1378_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1447_ _1441_/Y _1445_/Y _1446_/X VGND VGND VPWR VPWR _2217_/D sky130_fd_sc_hd__a21oi_4
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1301_ _1297_/X _1300_/X _1040_/X VGND VGND VPWR VPWR _1301_/Y sky130_fd_sc_hd__a21oi_4
X_1232_ _2083_/Q VGND VGND VPWR VPWR _1232_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1094_ _1076_/B _1090_/X _1093_/Y VGND VGND VPWR VPWR _1094_/Y sky130_fd_sc_hd__o21ai_4
X_1163_ _2084_/Q VGND VGND VPWR VPWR _1163_/Y sky130_fd_sc_hd__inv_2
X_1996_ SCSN_fromHost VGND VGND VPWR VPWR SCSN_toClient sky130_fd_sc_hd__buf_2
XFILLER_60_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1781_ _2120_/Q _1821_/B _1826_/A _1726_/A VGND VGND VPWR VPWR _1782_/A sky130_fd_sc_hd__and4_4
X_1850_ _1850_/A VGND VGND VPWR VPWR _1850_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1215_ _1215_/A _1215_/B _1190_/X VGND VGND VPWR VPWR _1215_/Y sky130_fd_sc_hd__nor3_4
X_1146_ _1182_/C VGND VGND VPWR VPWR _1215_/A sky130_fd_sc_hd__buf_2
XFILLER_37_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2195_ _2218_/CLK _2195_/D VGND VGND VPWR VPWR _1544_/A sky130_fd_sc_hd__dfxtp_4
X_1077_ _1059_/B _1076_/X _1072_/Y VGND VGND VPWR VPWR _1077_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1979_ PLL_INPUT M1_CLK_SELECT _1978_/Y VGND VGND VPWR VPWR m1_clk_local sky130_fd_sc_hd__o21a_4
XFILLER_20_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1000_ _1280_/A VGND VGND VPWR VPWR _1001_/A sky130_fd_sc_hd__buf_2
XFILLER_34_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1902_ _1902_/A VGND VGND VPWR VPWR _1902_/Y sky130_fd_sc_hd__inv_2
X_1833_ _2116_/Q _1832_/Y VGND VGND VPWR VPWR _1833_/Y sky130_fd_sc_hd__xnor2_4
X_1764_ _1746_/A _1762_/Y _1763_/Y VGND VGND VPWR VPWR _2134_/D sky130_fd_sc_hd__o21ai_4
X_1695_ _1694_/X _1695_/B VGND VGND VPWR VPWR _2154_/D sky130_fd_sc_hd__or2_4
X_1129_ _1108_/X _1087_/Y _1091_/X _1089_/X _1071_/X VGND VGND VPWR VPWR _1129_/Y
+ sky130_fd_sc_hd__a41oi_4
X_2247_ _2052_/CLK _2247_/D VGND VGND VPWR VPWR _2247_/Q sky130_fd_sc_hd__dfxtp_4
X_2178_ _2182_/CLK _2178_/D VGND VGND VPWR VPWR _1624_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_21_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9_0_addressalyzerBlock.SPI_CLK clkbuf_4_9_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2213_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1480_ _1480_/A _1480_/B VGND VGND VPWR VPWR _1480_/X sky130_fd_sc_hd__and2_4
X_2032_ _2124_/CLK _2038_/Q VGND VGND VPWR VPWR HASH_ADDR[1] sky130_fd_sc_hd__dfxtp_4
XFILLER_62_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2101_ _2108_/CLK _1862_/X VGND VGND VPWR VPWR _2101_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1816_ _1813_/A _1816_/B VGND VGND VPWR VPWR _2123_/D sky130_fd_sc_hd__xor2_4
X_1678_ _1678_/A _1668_/X VGND VGND VPWR VPWR _2164_/D sky130_fd_sc_hd__nor2_4
X_1747_ _1739_/X _1930_/A _1746_/Y VGND VGND VPWR VPWR _1747_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_42_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1601_ _1600_/Y VGND VGND VPWR VPWR _1601_/Y sky130_fd_sc_hd__inv_2
X_1532_ _2200_/Q _1525_/X _1531_/X VGND VGND VPWR VPWR _2201_/D sky130_fd_sc_hd__o21a_4
X_1394_ _1312_/X _1821_/B _1313_/B _1366_/A VGND VGND VPWR VPWR _1394_/X sky130_fd_sc_hd__a211o_4
X_1463_ _1412_/A _1462_/Y VGND VGND VPWR VPWR _1463_/Y sky130_fd_sc_hd__nor2_4
X_2015_ _2248_/CLK _1957_/Y VGND VGND VPWR VPWR _1451_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_23_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_1_0_m1_clk_local clkbuf_2_1_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_3_3_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_0_0_addressalyzerBlock.SPI_CLK clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_3_1_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
X_1515_ _1503_/X _1316_/A _1510_/X VGND VGND VPWR VPWR _1515_/X sky130_fd_sc_hd__o21a_4
X_1377_ _1153_/A VGND VGND VPWR VPWR _1473_/B sky130_fd_sc_hd__buf_2
X_1446_ _1098_/X VGND VGND VPWR VPWR _1446_/X sky130_fd_sc_hd__buf_2
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1300_ _1298_/Y _1299_/Y _1291_/X VGND VGND VPWR VPWR _1300_/X sky130_fd_sc_hd__a21o_4
X_1231_ _1159_/X _1484_/B _1161_/X VGND VGND VPWR VPWR _1231_/Y sky130_fd_sc_hd__a21oi_4
X_1162_ _1159_/X _1944_/C _1161_/X VGND VGND VPWR VPWR _1162_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_45_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1093_ _1076_/B _1053_/X _1091_/X _1090_/D _1957_/C VGND VGND VPWR VPWR _1093_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1995_ SCLK_fromHost VGND VGND VPWR VPWR SCLK_toClient sky130_fd_sc_hd__buf_2
X_1429_ _1427_/Y _1428_/X _1282_/C VGND VGND VPWR VPWR _1429_/X sky130_fd_sc_hd__o21a_4
XFILLER_55_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1780_ _1770_/Y _1780_/B _1840_/B VGND VGND VPWR VPWR _1825_/A sky130_fd_sc_hd__nor3_4
X_1145_ _1217_/A VGND VGND VPWR VPWR _1153_/A sky130_fd_sc_hd__inv_2
X_1214_ _1344_/C _1344_/D VGND VGND VPWR VPWR _1215_/B sky130_fd_sc_hd__nand2_4
XFILLER_37_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2194_ _2194_/CLK _2194_/D VGND VGND VPWR VPWR _1455_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1076_ _1053_/X _1076_/B _1125_/A _1090_/D VGND VGND VPWR VPWR _1076_/X sky130_fd_sc_hd__and4_4
XFILLER_33_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1978_ _1977_/Y M1_CLK_SELECT VGND VGND VPWR VPWR _1978_/Y sky130_fd_sc_hd__nand2_4
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1832_ _2115_/Q _1832_/B _1832_/C _1832_/D VGND VGND VPWR VPWR _1832_/Y sky130_fd_sc_hd__nand4_4
XFILLER_34_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1901_ _1316_/Y _1885_/X _1888_/X _1351_/Y _1890_/X VGND VGND VPWR VPWR _1901_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1763_ _1754_/A _1754_/B _1763_/C VGND VGND VPWR VPWR _1763_/Y sky130_fd_sc_hd__nand3_4
X_1694_ _1098_/A VGND VGND VPWR VPWR _1694_/X sky130_fd_sc_hd__buf_2
XFILLER_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2246_ _2052_/CLK _2246_/D VGND VGND VPWR VPWR _2246_/Q sky130_fd_sc_hd__dfxtp_4
X_1128_ _1128_/A _1069_/B VGND VGND VPWR VPWR _1128_/Y sky130_fd_sc_hd__nand2_4
X_1059_ _1090_/D _1059_/B _1076_/B _1105_/B VGND VGND VPWR VPWR _1059_/X sky130_fd_sc_hd__and4_4
X_2177_ _2171_/CLK _1635_/Y VGND VGND VPWR VPWR _1609_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_13_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_14_0_addressalyzerBlock.SPI_CLK clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2248_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_56_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2100_ _2091_/CLK _2100_/D VGND VGND VPWR VPWR _1867_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_62_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2031_ _2029_/CLK _2037_/Q VGND VGND VPWR VPWR HASH_ADDR[0] sky130_fd_sc_hd__dfxtp_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1815_ _1825_/A _1815_/B _1815_/C VGND VGND VPWR VPWR _1816_/B sky130_fd_sc_hd__and3_4
X_1677_ _1668_/X _1670_/B _1676_/Y VGND VGND VPWR VPWR _1677_/X sky130_fd_sc_hd__o21a_4
X_1746_ _1746_/A _1969_/A _1230_/A VGND VGND VPWR VPWR _1746_/Y sky130_fd_sc_hd__nand3_4
X_2229_ _2058_/CLK _1287_/Y VGND VGND VPWR VPWR _1178_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_53_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1600_ _1589_/B _1600_/B _1600_/C VGND VGND VPWR VPWR _1600_/Y sky130_fd_sc_hd__nand3_4
XFILLER_4_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1531_ _2201_/Q _1526_/X _1521_/X VGND VGND VPWR VPWR _1531_/X sky130_fd_sc_hd__o21a_4
XFILLER_8_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1462_ _1462_/A VGND VGND VPWR VPWR _1462_/Y sky130_fd_sc_hd__inv_2
X_1393_ _1391_/Y _1285_/X _1392_/Y VGND VGND VPWR VPWR _1393_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_50_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2014_ _2248_/CLK _1965_/Y VGND VGND VPWR VPWR _2014_/Q sky130_fd_sc_hd__dfxtp_4
X_1729_ _1310_/A _1847_/A _1202_/Y _1243_/B _1270_/Y VGND VGND VPWR VPWR _1729_/Y
+ sky130_fd_sc_hd__o41ai_4
XFILLER_58_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1445_ _1445_/A _1957_/B _1444_/Y _1449_/C VGND VGND VPWR VPWR _1445_/Y sky130_fd_sc_hd__nand4_4
X_1514_ _1573_/B _2200_/Q _1513_/X VGND VGND VPWR VPWR _2208_/D sky130_fd_sc_hd__o21a_4
XFILLER_55_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1376_ _1376_/A VGND VGND VPWR VPWR _1788_/A sky130_fd_sc_hd__inv_2
XFILLER_23_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1092_ _1092_/A VGND VGND VPWR VPWR _1957_/C sky130_fd_sc_hd__buf_2
X_1230_ _1230_/A _1155_/X VGND VGND VPWR VPWR _1230_/Y sky130_fd_sc_hd__nand2_4
X_1161_ _1161_/A VGND VGND VPWR VPWR _1161_/X sky130_fd_sc_hd__buf_2
X_1994_ MOSI_fromHost VGND VGND VPWR VPWR MOSI_toClient sky130_fd_sc_hd__buf_2
XFILLER_20_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1428_ _1001_/A _1972_/C VGND VGND VPWR VPWR _1428_/X sky130_fd_sc_hd__or2_4
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1359_ _1354_/X _1358_/X VGND VGND VPWR VPWR _1359_/Y sky130_fd_sc_hd__nand2_4
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1213_ _1213_/A VGND VGND VPWR VPWR _1226_/A sky130_fd_sc_hd__inv_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1144_ _1311_/A _1144_/B VGND VGND VPWR VPWR _1217_/A sky130_fd_sc_hd__nor2_4
X_1075_ _1105_/B VGND VGND VPWR VPWR _1125_/A sky130_fd_sc_hd__buf_2
XFILLER_37_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2193_ _2194_/CLK _2193_/D VGND VGND VPWR VPWR _1455_/D sky130_fd_sc_hd__dfxtp_4
X_1977_ M1_CLK_IN VGND VGND VPWR VPWR _1977_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1831_ _1770_/Y VGND VGND VPWR VPWR _1832_/D sky130_fd_sc_hd__inv_2
XFILLER_42_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1900_ _1112_/Y _1899_/A _1899_/Y VGND VGND VPWR VPWR _1900_/Y sky130_fd_sc_hd__o21ai_4
X_1762_ _1504_/X _1445_/A _1133_/X VGND VGND VPWR VPWR _1762_/Y sky130_fd_sc_hd__nand3_4
X_1693_ _1704_/A _1693_/B _1702_/B _1693_/D VGND VGND VPWR VPWR _1693_/X sky130_fd_sc_hd__and4_4
X_2245_ _2052_/CLK _1019_/Y VGND VGND VPWR VPWR _2245_/Q sky130_fd_sc_hd__dfxtp_4
X_2176_ _2171_/CLK _2176_/D VGND VGND VPWR VPWR _1576_/A sky130_fd_sc_hd__dfxtp_4
X_1127_ _1326_/A _1123_/X _1126_/Y VGND VGND VPWR VPWR _1128_/A sky130_fd_sc_hd__a21o_4
X_1058_ _1097_/A VGND VGND VPWR VPWR _1076_/B sky130_fd_sc_hd__buf_2
XFILLER_25_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2030_ _2029_/CLK _2030_/D VGND VGND VPWR VPWR _2029_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_62_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1814_ _2124_/Q _1813_/Y VGND VGND VPWR VPWR _1814_/Y sky130_fd_sc_hd__xnor2_4
X_1745_ _1633_/A _1740_/X _1892_/A VGND VGND VPWR VPWR _1930_/A sky130_fd_sc_hd__nand3_4
X_1676_ _1668_/X _1670_/B _1102_/A VGND VGND VPWR VPWR _1676_/Y sky130_fd_sc_hd__a21oi_4
X_2228_ _2228_/CLK _2228_/D VGND VGND VPWR VPWR _1147_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_26_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2159_ _2194_/CLK _1686_/X VGND VGND VPWR VPWR _1983_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_53_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_0_0_addressalyzerBlock.SPI_CLK clkbuf_3_1_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_4_1_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_13_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1392_ _1179_/X _2047_/Q _1188_/X VGND VGND VPWR VPWR _1392_/Y sky130_fd_sc_hd__o21ai_4
X_1461_ _1459_/Y _1460_/Y _1052_/B VGND VGND VPWR VPWR _1461_/X sky130_fd_sc_hd__a21o_4
X_1530_ _2201_/Q _1525_/X _1529_/X VGND VGND VPWR VPWR _1530_/X sky130_fd_sc_hd__o21a_4
X_2013_ _2248_/CLK _1968_/X VGND VGND VPWR VPWR _1451_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_35_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1728_ _2109_/Q VGND VGND VPWR VPWR _1847_/A sky130_fd_sc_hd__inv_2
X_1659_ _1659_/A VGND VGND VPWR VPWR _1659_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1375_ _1343_/X _1373_/Y _1374_/Y VGND VGND VPWR VPWR _1375_/Y sky130_fd_sc_hd__o21ai_4
X_1444_ _1451_/B VGND VGND VPWR VPWR _1444_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1513_ _1503_/X _1112_/A _1510_/X VGND VGND VPWR VPWR _1513_/X sky130_fd_sc_hd__o21a_4
XFILLER_23_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1091_ _1125_/A VGND VGND VPWR VPWR _1091_/X sky130_fd_sc_hd__buf_2
XFILLER_38_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1160_ _2144_/Q VGND VGND VPWR VPWR _1161_/A sky130_fd_sc_hd__inv_2
XFILLER_60_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1993_ EXT_RESET_N_fromHost VGND VGND VPWR VPWR EXT_RESET_N_toClient sky130_fd_sc_hd__buf_2
XFILLER_9_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1427_ _1308_/X _1431_/A VGND VGND VPWR VPWR _1427_/Y sky130_fd_sc_hd__nor2_4
X_1358_ _1757_/C _1155_/X _1161_/X _1357_/Y VGND VGND VPWR VPWR _1358_/X sky130_fd_sc_hd__a211o_4
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1289_ _1125_/D _1105_/A _1288_/X VGND VGND VPWR VPWR _1289_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_36_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2192_ _2189_/CLK _2192_/D VGND VGND VPWR VPWR _2192_/Q sky130_fd_sc_hd__dfxtp_4
X_1212_ _1834_/B VGND VGND VPWR VPWR _1212_/Y sky130_fd_sc_hd__inv_2
X_1143_ _1048_/D VGND VGND VPWR VPWR _1144_/B sky130_fd_sc_hd__inv_2
X_1074_ _1069_/Y _1073_/Y _1040_/X VGND VGND VPWR VPWR _2240_/D sky130_fd_sc_hd__a21oi_4
XFILLER_33_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1976_ EXT_RESET_N_fromHost VGND VGND VPWR VPWR _1976_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1830_ _1829_/X VGND VGND VPWR VPWR _1832_/B sky130_fd_sc_hd__buf_2
XFILLER_30_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1761_ _1746_/A _1759_/Y _1760_/Y VGND VGND VPWR VPWR _1761_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_15_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1692_ _1692_/A VGND VGND VPWR VPWR _1702_/B sky130_fd_sc_hd__inv_2
X_2244_ _2052_/CLK _2244_/D VGND VGND VPWR VPWR _1020_/A sky130_fd_sc_hd__dfxtp_4
X_2175_ _2182_/CLK _1640_/Y VGND VGND VPWR VPWR _2175_/Q sky130_fd_sc_hd__dfxtp_4
X_1126_ _1116_/B _1126_/B _1071_/X _1126_/D VGND VGND VPWR VPWR _1126_/Y sky130_fd_sc_hd__nor4_4
X_1057_ _1057_/A _2236_/Q _2235_/Q _1108_/A VGND VGND VPWR VPWR _1090_/D sky130_fd_sc_hd__and4_4
XFILLER_25_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1959_ _1694_/X _1036_/B _1972_/C _1971_/C _1958_/Y VGND VGND VPWR VPWR _1959_/Y
+ sky130_fd_sc_hd__o41ai_4
XFILLER_48_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_6_0_m1_clk_local clkbuf_3_7_0_m1_clk_local/A VGND VGND VPWR VPWR _2025_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1813_ _1813_/A _1827_/B _1815_/B _1815_/C VGND VGND VPWR VPWR _1813_/Y sky130_fd_sc_hd__nand4_4
XFILLER_7_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1744_ _1739_/X _1741_/Y _1743_/Y VGND VGND VPWR VPWR _2140_/D sky130_fd_sc_hd__o21ai_4
X_1675_ _1674_/X _1675_/B _1675_/C VGND VGND VPWR VPWR _2166_/D sky130_fd_sc_hd__and3_4
X_2227_ _2216_/CLK _1301_/Y VGND VGND VPWR VPWR _1149_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1109_ _1109_/A _1106_/X _1116_/B _1108_/X VGND VGND VPWR VPWR _1109_/Y sky130_fd_sc_hd__nand4_4
X_2089_ _2213_/CLK _1900_/Y VGND VGND VPWR VPWR _2001_/D sky130_fd_sc_hd__dfxtp_4
X_2158_ _2218_/CLK _1689_/X VGND VGND VPWR VPWR _2158_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1391_ _1386_/X _1390_/X VGND VGND VPWR VPWR _1391_/Y sky130_fd_sc_hd__nand2_4
X_1460_ _1460_/A _1355_/X VGND VGND VPWR VPWR _1460_/Y sky130_fd_sc_hd__nand2_4
X_2012_ _2248_/CLK _2012_/D VGND VGND VPWR VPWR _2012_/Q sky130_fd_sc_hd__dfxtp_4
X_1727_ _1312_/X _1825_/B _1313_/B _1362_/A VGND VGND VPWR VPWR _1727_/X sky130_fd_sc_hd__a211o_4
X_1658_ _1648_/X _1649_/A _1657_/Y VGND VGND VPWR VPWR _1659_/A sky130_fd_sc_hd__o21ai_4
XFILLER_58_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1589_ _1589_/A _1589_/B _1589_/C _2185_/Q VGND VGND VPWR VPWR _1589_/Y sky130_fd_sc_hd__nand4_4
XFILLER_53_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1512_ _1573_/B _2201_/Q _1511_/X VGND VGND VPWR VPWR _1512_/X sky130_fd_sc_hd__o21a_4
XFILLER_55_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1374_ _1274_/A _1374_/B VGND VGND VPWR VPWR _1374_/Y sky130_fd_sc_hd__nand2_4
X_1443_ _1442_/X VGND VGND VPWR VPWR _1445_/A sky130_fd_sc_hd__buf_2
XFILLER_23_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1090_ _1087_/Y _1125_/A _1089_/X _1090_/D VGND VGND VPWR VPWR _1090_/X sky130_fd_sc_hd__and4_4
X_1992_ VGND VGND VPWR VPWR _1992_/HI zero sky130_fd_sc_hd__conb_1
XFILLER_20_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1288_ _1084_/Y _1085_/Y _1086_/X _1049_/X _1298_/C VGND VGND VPWR VPWR _1288_/X
+ sky130_fd_sc_hd__o41a_4
X_1357_ _1355_/X _1356_/Y VGND VGND VPWR VPWR _1357_/Y sky130_fd_sc_hd__nor2_4
X_1426_ _1426_/A VGND VGND VPWR VPWR _1426_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2191_ _2189_/CLK _2191_/D VGND VGND VPWR VPWR _1563_/A sky130_fd_sc_hd__dfxtp_4
X_1211_ _1779_/A VGND VGND VPWR VPWR _1834_/B sky130_fd_sc_hd__buf_2
X_1142_ _1138_/Y _1140_/Y _1141_/Y VGND VGND VPWR VPWR _1142_/Y sky130_fd_sc_hd__a21oi_4
X_1073_ _1070_/X _1072_/Y _2240_/Q VGND VGND VPWR VPWR _1073_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_33_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1975_ _1974_/X _1436_/Y _1701_/A VGND VGND VPWR VPWR _1975_/X sky130_fd_sc_hd__o21a_4
X_1409_ _1407_/Y _1233_/X _1408_/Y VGND VGND VPWR VPWR _1409_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_43_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_0_0_addressalyzerBlock.SPI_CLK clkbuf_4_1_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2091_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_15_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1760_ _1754_/A _1754_/B _1760_/C VGND VGND VPWR VPWR _1760_/Y sky130_fd_sc_hd__nand3_4
X_1691_ _1656_/A _1692_/A _1693_/D _1693_/B VGND VGND VPWR VPWR _2156_/D sky130_fd_sc_hd__nor4_4
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1125_ _1125_/A _1105_/A _1088_/X _1125_/D VGND VGND VPWR VPWR _1126_/D sky130_fd_sc_hd__nand4_4
X_2243_ _2052_/CLK _1027_/Y VGND VGND VPWR VPWR _1024_/A sky130_fd_sc_hd__dfxtp_4
X_2174_ _2182_/CLK _2174_/D VGND VGND VPWR VPWR _2174_/Q sky130_fd_sc_hd__dfxtp_4
X_1056_ _1092_/A VGND VGND VPWR VPWR _1110_/A sky130_fd_sc_hd__inv_2
XFILLER_21_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1958_ _1958_/A _1044_/Y _1001_/A _1969_/D VGND VGND VPWR VPWR _1958_/Y sky130_fd_sc_hd__nand4_4
X_1889_ _1329_/X _1219_/B _1195_/X _1442_/X _1330_/A VGND VGND VPWR VPWR _1889_/X
+ sky130_fd_sc_hd__a41o_4
Xclkbuf_3_5_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1812_ _1825_/A VGND VGND VPWR VPWR _1827_/B sky130_fd_sc_hd__buf_2
X_1674_ _1668_/A _1670_/B _2166_/Q VGND VGND VPWR VPWR _1674_/X sky130_fd_sc_hd__a21o_4
X_1743_ _1746_/A _1969_/A _1156_/A VGND VGND VPWR VPWR _1743_/Y sky130_fd_sc_hd__nand3_4
X_2226_ _2231_/CLK _1307_/X VGND VGND VPWR VPWR _1149_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_53_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1108_ _1108_/A VGND VGND VPWR VPWR _1108_/X sky130_fd_sc_hd__buf_2
X_1039_ _1098_/A VGND VGND VPWR VPWR _1040_/A sky130_fd_sc_hd__buf_2
X_2157_ _2248_/CLK _1690_/Y VGND VGND VPWR VPWR _1972_/C sky130_fd_sc_hd__dfxtp_4
X_2088_ _2085_/CLK _1901_/Y VGND VGND VPWR VPWR _2088_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_29_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1390_ _1760_/C _1155_/X _1161_/A _1389_/Y VGND VGND VPWR VPWR _1390_/X sky130_fd_sc_hd__a211o_4
XFILLER_50_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2011_ _2216_/CLK _2011_/D VGND VGND VPWR VPWR _1064_/A sky130_fd_sc_hd__dfxtp_4
X_1726_ _1726_/A VGND VGND VPWR VPWR _1825_/B sky130_fd_sc_hd__buf_2
X_1657_ _1649_/A _1648_/X _1293_/X VGND VGND VPWR VPWR _1657_/Y sky130_fd_sc_hd__a21oi_4
X_1588_ _1595_/A _1588_/B VGND VGND VPWR VPWR _1589_/B sky130_fd_sc_hd__nor2_4
XFILLER_58_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2209_ _2211_/CLK _1512_/X VGND VGND VPWR VPWR _1748_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1511_ _1503_/X _1894_/A _1510_/X VGND VGND VPWR VPWR _1511_/X sky130_fd_sc_hd__o21a_4
X_1442_ _2217_/Q VGND VGND VPWR VPWR _1442_/X sky130_fd_sc_hd__buf_2
X_1373_ THREAD_COUNT[3] _1421_/A _1369_/Y _1372_/Y VGND VGND VPWR VPWR _1373_/Y sky130_fd_sc_hd__a22oi_4
X_1709_ _1217_/X _1708_/A _1215_/Y _1708_/X VGND VGND VPWR VPWR _1709_/X sky130_fd_sc_hd__a211o_4
XFILLER_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1991_ VGND VGND VPWR VPWR one _1991_/LO sky130_fd_sc_hd__conb_1
X_1425_ _1343_/X _1423_/Y _1424_/Y VGND VGND VPWR VPWR _2219_/D sky130_fd_sc_hd__o21ai_4
X_1287_ _1277_/Y _1284_/Y _1286_/X VGND VGND VPWR VPWR _1287_/Y sky130_fd_sc_hd__a21oi_4
X_1356_ _2064_/Q VGND VGND VPWR VPWR _1356_/Y sky130_fd_sc_hd__inv_2
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2190_ _2189_/CLK _1568_/X VGND VGND VPWR VPWR _1562_/C sky130_fd_sc_hd__dfxtp_4
X_1210_ _1203_/Y _2116_/Q _1209_/X VGND VGND VPWR VPWR _1210_/Y sky130_fd_sc_hd__a21oi_4
X_1141_ _1091_/X _1069_/B _1031_/X VGND VGND VPWR VPWR _1141_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_37_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1072_ _1053_/X _1061_/D _1071_/X VGND VGND VPWR VPWR _1072_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_60_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1974_ _1308_/X _1451_/A _1451_/C VGND VGND VPWR VPWR _1974_/X sky130_fd_sc_hd__o21a_4
X_1408_ _1171_/X _2038_/D _1172_/X VGND VGND VPWR VPWR _1408_/Y sky130_fd_sc_hd__a21oi_4
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1339_ _1291_/X _1144_/B VGND VGND VPWR VPWR _1341_/B sky130_fd_sc_hd__nand2_4
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1690_ _1656_/A _2148_/Q _1688_/Y VGND VGND VPWR VPWR _1690_/Y sky130_fd_sc_hd__nor3_4
X_2242_ _2052_/CLK _1033_/Y VGND VGND VPWR VPWR _2242_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2173_ _2189_/CLK _1651_/X VGND VGND VPWR VPWR _2173_/Q sky130_fd_sc_hd__dfxtp_4
X_1055_ _1055_/A VGND VGND VPWR VPWR _1092_/A sky130_fd_sc_hd__buf_2
X_1124_ _1108_/A VGND VGND VPWR VPWR _1126_/B sky130_fd_sc_hd__inv_2
X_1957_ _1656_/A _1957_/B _1957_/C VGND VGND VPWR VPWR _1957_/Y sky130_fd_sc_hd__nor3_4
X_1888_ _1887_/Y VGND VGND VPWR VPWR _1888_/X sky130_fd_sc_hd__buf_2
XFILLER_56_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1811_ _1803_/A _1787_/Y VGND VGND VPWR VPWR _2125_/D sky130_fd_sc_hd__xor2_4
XFILLER_30_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1673_ _2167_/Q _1671_/Y _1672_/Y VGND VGND VPWR VPWR _1673_/X sky130_fd_sc_hd__o21a_4
X_1742_ _1738_/Y VGND VGND VPWR VPWR _1746_/A sky130_fd_sc_hd__buf_2
XFILLER_7_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2225_ _2231_/CLK _1324_/Y VGND VGND VPWR VPWR _1182_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_53_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1107_ _2235_/Q VGND VGND VPWR VPWR _1116_/B sky130_fd_sc_hd__buf_2
X_2087_ _2091_/CLK _2087_/D VGND VGND VPWR VPWR _1383_/A sky130_fd_sc_hd__dfxtp_4
X_2156_ _2194_/CLK _2156_/D VGND VGND VPWR VPWR _2156_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_21_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1038_ _1038_/A VGND VGND VPWR VPWR _1098_/A sky130_fd_sc_hd__buf_2
XFILLER_44_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2010_ _2216_/CLK _1970_/Y VGND VGND VPWR VPWR _2010_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_3_2_0_m1_clk_local clkbuf_3_3_0_m1_clk_local/A VGND VGND VPWR VPWR _2189_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_1725_ _1711_/Y _1723_/Y _1724_/Y VGND VGND VPWR VPWR _1725_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_58_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1656_ _1656_/A _1583_/B _1656_/C VGND VGND VPWR VPWR _2171_/D sky130_fd_sc_hd__nor3_4
X_1587_ _1587_/A _1584_/Y _2181_/Q _1587_/D VGND VGND VPWR VPWR _1588_/B sky130_fd_sc_hd__nand4_4
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2139_ _2137_/CLK _1747_/Y VGND VGND VPWR VPWR _1230_/A sky130_fd_sc_hd__dfxtp_4
X_2208_ _2211_/CLK _2208_/D VGND VGND VPWR VPWR _1112_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_26_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1510_ _1633_/A VGND VGND VPWR VPWR _1510_/X sky130_fd_sc_hd__buf_2
X_1441_ _1436_/Y _1438_/Y _1440_/X VGND VGND VPWR VPWR _1441_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_63_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1372_ _1209_/X _1371_/X _1421_/A VGND VGND VPWR VPWR _1372_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_48_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1708_ _1708_/A THREAD_COUNT[0] _1344_/A VGND VGND VPWR VPWR _1708_/X sky130_fd_sc_hd__and3_4
X_1639_ _1607_/X _1646_/C _1031_/X VGND VGND VPWR VPWR _1639_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1990_ _1988_/Y _1030_/X _1989_/Y VGND VGND VPWR VPWR _1990_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1424_ _1480_/A _2219_/Q VGND VGND VPWR VPWR _1424_/Y sky130_fd_sc_hd__nand2_4
X_1355_ _1355_/A VGND VGND VPWR VPWR _1355_/X sky130_fd_sc_hd__buf_2
XFILLER_55_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1286_ _1306_/A _1285_/X _1098_/X VGND VGND VPWR VPWR _1286_/X sky130_fd_sc_hd__a21o_4
XFILLER_36_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_5_0_addressalyzerBlock.SPI_CLK clkbuf_4_5_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2044_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_52_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1071_ _1092_/A VGND VGND VPWR VPWR _1071_/X sky130_fd_sc_hd__buf_2
X_1140_ _1907_/A _1123_/X _1079_/X VGND VGND VPWR VPWR _1140_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_60_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1973_ _1553_/Y _1065_/A _1694_/X _1972_/X VGND VGND VPWR VPWR _1973_/X sky130_fd_sc_hd__a211o_4
X_1338_ _1907_/A _1279_/Y _1337_/X _1291_/A VGND VGND VPWR VPWR _1341_/A sky130_fd_sc_hd__a211o_4
X_1407_ _1998_/D VGND VGND VPWR VPWR _1407_/Y sky130_fd_sc_hd__inv_2
X_1269_ _1203_/Y _1770_/A _1209_/X VGND VGND VPWR VPWR _1269_/Y sky130_fd_sc_hd__a21oi_4
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2241_ _2052_/CLK _1041_/Y VGND VGND VPWR VPWR _1034_/C sky130_fd_sc_hd__dfxtp_4
X_2172_ _2171_/CLK _2172_/D VGND VGND VPWR VPWR _1583_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_33_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1054_ _2010_/Q _1449_/B VGND VGND VPWR VPWR _1055_/A sky130_fd_sc_hd__nor2_4
X_1123_ _2012_/Q VGND VGND VPWR VPWR _1123_/X sky130_fd_sc_hd__buf_2
XFILLER_25_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1887_ _1887_/A VGND VGND VPWR VPWR _1887_/Y sky130_fd_sc_hd__inv_2
X_1956_ _1719_/Y _1948_/X _1907_/A _1943_/A VGND VGND VPWR VPWR _1956_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1810_ _1810_/A _1810_/B VGND VGND VPWR VPWR _2126_/D sky130_fd_sc_hd__xor2_4
X_1741_ _1917_/A _1740_/X _1042_/A VGND VGND VPWR VPWR _1741_/Y sky130_fd_sc_hd__nand3_4
X_1672_ _1668_/X _1670_/B _2166_/Q _2167_/Q _1040_/A VGND VGND VPWR VPWR _1672_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1106_ _1106_/A VGND VGND VPWR VPWR _1106_/X sky130_fd_sc_hd__buf_2
XFILLER_26_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2224_ _2224_/CLK _2224_/D VGND VGND VPWR VPWR _1184_/A sky130_fd_sc_hd__dfxtp_4
X_2155_ _2218_/CLK _1693_/X VGND VGND VPWR VPWR _0995_/A sky130_fd_sc_hd__dfxtp_4
X_2086_ _2085_/CLK _2086_/D VGND VGND VPWR VPWR _1998_/D sky130_fd_sc_hd__dfxtp_4
X_1037_ _2006_/Q VGND VGND VPWR VPWR _1038_/A sky130_fd_sc_hd__buf_2
X_1939_ _1904_/Y _1934_/Y _1733_/D _1404_/Y _1935_/Y VGND VGND VPWR VPWR _2070_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0_addressalyzerBlock.SPI_CLK clkbuf_0_addressalyzerBlock.SPI_CLK/X VGND
+ VGND VPWR VPWR clkbuf_2_3_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_4_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1724_ _1186_/Y _1769_/A _1153_/Y VGND VGND VPWR VPWR _1724_/Y sky130_fd_sc_hd__a21oi_4
X_1655_ _1649_/A _1648_/X _1649_/C VGND VGND VPWR VPWR _1656_/C sky130_fd_sc_hd__a21oi_4
X_1586_ _1585_/Y VGND VGND VPWR VPWR _1587_/D sky130_fd_sc_hd__inv_2
X_2138_ _2137_/CLK _1752_/Y VGND VGND VPWR VPWR _1253_/A sky130_fd_sc_hd__dfxtp_4
X_2069_ _2211_/CLK _1941_/X VGND VGND VPWR VPWR _2030_/D sky130_fd_sc_hd__dfxtp_4
X_2207_ _2211_/CLK _1516_/X VGND VGND VPWR VPWR _1316_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_34_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1371_ _1371_/A VGND VGND VPWR VPWR _1371_/X sky130_fd_sc_hd__buf_2
X_1440_ _1886_/C _1298_/C _2213_/Q _1451_/A VGND VGND VPWR VPWR _1440_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1707_ _1341_/Y VGND VGND VPWR VPWR _2142_/D sky130_fd_sc_hd__inv_2
X_1638_ _1637_/Y VGND VGND VPWR VPWR _2176_/D sky130_fd_sc_hd__inv_2
X_1569_ _1569_/A _2189_/Q VGND VGND VPWR VPWR _1569_/X sky130_fd_sc_hd__or2_4
XFILLER_39_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1423_ THREAD_COUNT[1] _1421_/A _1420_/Y _1422_/X VGND VGND VPWR VPWR _1423_/Y sky130_fd_sc_hd__a22oi_4
X_1285_ _1178_/Y VGND VGND VPWR VPWR _1285_/X sky130_fd_sc_hd__buf_2
X_1354_ _1350_/X _1353_/Y _1175_/X VGND VGND VPWR VPWR _1354_/X sky130_fd_sc_hd__a21o_4
XFILLER_27_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_10_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2194_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_54_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1070_ _1067_/Y VGND VGND VPWR VPWR _1070_/X sky130_fd_sc_hd__buf_2
XFILLER_1_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1972_ _1972_/A _1004_/A _1972_/C VGND VGND VPWR VPWR _1972_/X sky130_fd_sc_hd__and3_4
X_1268_ _1153_/Y _1266_/Y _1267_/X VGND VGND VPWR VPWR _1268_/Y sky130_fd_sc_hd__o21ai_4
X_1337_ _2010_/Q _1449_/B _1144_/B VGND VGND VPWR VPWR _1337_/X sky130_fd_sc_hd__o21a_4
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1406_ _2078_/Q _1154_/X _1166_/X _1405_/Y VGND VGND VPWR VPWR _1406_/X sky130_fd_sc_hd__a211o_4
XFILLER_61_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1199_ _1195_/X _2124_/Q _1196_/X _1473_/C VGND VGND VPWR VPWR _1199_/X sky130_fd_sc_hd__a211o_4
XFILLER_51_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2171_ _2171_/CLK _2171_/D VGND VGND VPWR VPWR _1643_/A sky130_fd_sc_hd__dfxtp_4
X_2240_ _2228_/CLK _2240_/D VGND VGND VPWR VPWR _2240_/Q sky130_fd_sc_hd__dfxtp_4
X_1122_ _1118_/Y _1119_/Y _1121_/X VGND VGND VPWR VPWR _1122_/Y sky130_fd_sc_hd__a21oi_4
X_1053_ _1052_/X VGND VGND VPWR VPWR _1053_/X sky130_fd_sc_hd__buf_2
XFILLER_33_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1955_ _1411_/Y _1949_/X _1133_/X _1950_/X VGND VGND VPWR VPWR _1955_/X sky130_fd_sc_hd__a2bb2o_4
X_1886_ _1038_/A _1310_/X _1886_/C VGND VGND VPWR VPWR _1887_/A sky130_fd_sc_hd__nor3_4
XFILLER_56_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1671_ _1675_/C VGND VGND VPWR VPWR _1671_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1740_ _1442_/X VGND VGND VPWR VPWR _1740_/X sky130_fd_sc_hd__buf_2
XFILLER_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1105_ _1105_/A _1105_/B _1178_/A _1147_/B VGND VGND VPWR VPWR _1106_/A sky130_fd_sc_hd__and4_4
XFILLER_38_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2223_ _2216_/CLK _2223_/D VGND VGND VPWR VPWR _1047_/A sky130_fd_sc_hd__dfxtp_4
X_2085_ _2085_/CLK _1908_/Y VGND VGND VPWR VPWR _1997_/D sky130_fd_sc_hd__dfxtp_4
X_2154_ _2218_/CLK _2154_/D VGND VGND VPWR VPWR _1692_/A sky130_fd_sc_hd__dfxtp_4
X_1036_ _2141_/Q _1036_/B VGND VGND VPWR VPWR _1036_/Y sky130_fd_sc_hd__nand2_4
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1869_ _1867_/A _1767_/B _1869_/C VGND VGND VPWR VPWR _1869_/Y sky130_fd_sc_hd__nand3_4
X_1938_ _1902_/Y _1934_/Y _1733_/D _1380_/Y _1935_/Y VGND VGND VPWR VPWR _1938_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1723_ _1052_/B _1722_/Y VGND VGND VPWR VPWR _1723_/Y sky130_fd_sc_hd__nor2_4
X_1654_ _1330_/X VGND VGND VPWR VPWR _1656_/A sky130_fd_sc_hd__buf_2
X_2206_ _2194_/CLK _1518_/X VGND VGND VPWR VPWR _1326_/A sky130_fd_sc_hd__dfxtp_4
X_1585_ _1624_/D _1627_/D VGND VGND VPWR VPWR _1585_/Y sky130_fd_sc_hd__nand2_4
X_1019_ _1017_/Y _1003_/X _1018_/Y VGND VGND VPWR VPWR _1019_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_34_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2137_ _2137_/CLK _1755_/Y VGND VGND VPWR VPWR _1460_/A sky130_fd_sc_hd__dfxtp_4
X_2068_ _2085_/CLK _2068_/D VGND VGND VPWR VPWR _1944_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_57_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1370_ _1370_/A VGND VGND VPWR VPWR _1371_/A sky130_fd_sc_hd__inv_2
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1706_ _1318_/X _1323_/C _1333_/Y _1334_/Y _1335_/X VGND VGND VPWR VPWR _2143_/D
+ sky130_fd_sc_hd__a41oi_4
X_1637_ _1621_/B _1619_/Y _1636_/Y VGND VGND VPWR VPWR _1637_/Y sky130_fd_sc_hd__o21ai_4
X_1568_ _1570_/A SPI_CLK_RESET_N _1562_/Y _1568_/D VGND VGND VPWR VPWR _1568_/X sky130_fd_sc_hd__and4_4
X_1499_ _1426_/Y _1499_/B VGND VGND VPWR VPWR _1499_/Y sky130_fd_sc_hd__nand2_4
XFILLER_54_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1422_ _2102_/Q _1270_/Y _1421_/Y VGND VGND VPWR VPWR _1422_/X sky130_fd_sc_hd__o21a_4
X_1284_ _1042_/A _1279_/Y _1306_/A VGND VGND VPWR VPWR _1284_/Y sky130_fd_sc_hd__a21oi_4
X_1353_ _1351_/Y _1233_/X _1352_/Y VGND VGND VPWR VPWR _1353_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_63_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0999_ _2246_/Q _0996_/X _0998_/X VGND VGND VPWR VPWR _0999_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1971_ _1971_/A _1971_/B _1971_/C VGND VGND VPWR VPWR _1972_/A sky130_fd_sc_hd__nand3_4
XFILLER_5_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1405_ _1355_/A _1404_/Y VGND VGND VPWR VPWR _1405_/Y sky130_fd_sc_hd__nor2_4
X_1198_ _1362_/A VGND VGND VPWR VPWR _1473_/C sky130_fd_sc_hd__buf_2
X_1267_ _1195_/X _2122_/Q _1196_/X _1473_/C VGND VGND VPWR VPWR _1267_/X sky130_fd_sc_hd__a211o_4
X_1336_ _1318_/X _1323_/C _1333_/Y _1334_/Y _1335_/X VGND VGND VPWR VPWR _2223_/D
+ sky130_fd_sc_hd__a41oi_4
XFILLER_51_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_addressalyzerBlock.SPI_CLK _1982_/Y VGND VGND VPWR VPWR clkbuf_0_addressalyzerBlock.SPI_CLK/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_19_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1052_ _1052_/A _1052_/B _1147_/B _1149_/A VGND VGND VPWR VPWR _1052_/X sky130_fd_sc_hd__and4_4
X_2170_ _2124_/CLK _1659_/Y VGND VGND VPWR VPWR _1648_/A sky130_fd_sc_hd__dfxtp_4
X_1121_ _1070_/X _1120_/Y _1098_/X VGND VGND VPWR VPWR _1121_/X sky130_fd_sc_hd__a21o_4
XFILLER_33_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1954_ _1389_/B _1949_/X _1902_/A _1950_/X VGND VGND VPWR VPWR _1954_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_2_1_0_addressalyzerBlock.SPI_CLK clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
X_1885_ _1473_/B VGND VGND VPWR VPWR _1885_/X sky130_fd_sc_hd__buf_2
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1319_ _2010_/Q VGND VGND VPWR VPWR _1971_/A sky130_fd_sc_hd__inv_2
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1670_ _1668_/X _1670_/B _2166_/Q VGND VGND VPWR VPWR _1675_/C sky130_fd_sc_hd__nand3_4
X_2222_ _2228_/CLK _1342_/Y VGND VGND VPWR VPWR _1048_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1104_ _1085_/Y _1086_/A _1049_/A VGND VGND VPWR VPWR _1105_/A sky130_fd_sc_hd__nor3_4
XFILLER_38_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1035_ _1001_/A VGND VGND VPWR VPWR _1036_/B sky130_fd_sc_hd__buf_2
X_2153_ _2218_/CLK _1696_/X VGND VGND VPWR VPWR _1695_/B sky130_fd_sc_hd__dfxtp_4
X_2084_ _2085_/CLK _2084_/D VGND VGND VPWR VPWR _2084_/Q sky130_fd_sc_hd__dfxtp_4
X_1937_ _1316_/Y _1934_/Y _1733_/D _1348_/Y _1935_/Y VGND VGND VPWR VPWR _2072_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1799_ _1798_/X _1799_/B VGND VGND VPWR VPWR _1800_/A sky130_fd_sc_hd__nand2_4
X_1868_ _1741_/Y _1865_/X _1867_/Y VGND VGND VPWR VPWR _2100_/D sky130_fd_sc_hd__o21ai_4
XFILLER_16_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1653_ _1649_/D _1583_/B _1652_/Y VGND VGND VPWR VPWR _2172_/D sky130_fd_sc_hd__o21a_4
X_1584_ _1575_/Y _1584_/B _1584_/C _1583_/Y VGND VGND VPWR VPWR _1584_/Y sky130_fd_sc_hd__nor4_4
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1722_ _1718_/Y _1161_/X _1721_/X VGND VGND VPWR VPWR _1722_/Y sky130_fd_sc_hd__a21boi_4
X_2205_ _2213_/CLK _2205_/D VGND VGND VPWR VPWR _1904_/A sky130_fd_sc_hd__dfxtp_4
X_1018_ _1480_/B _1004_/X _1008_/X VGND VGND VPWR VPWR _1018_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_41_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2136_ _2137_/CLK _2136_/D VGND VGND VPWR VPWR _1757_/C sky130_fd_sc_hd__dfxtp_4
X_2067_ _2085_/CLK _2067_/D VGND VGND VPWR VPWR _1484_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1705_ _1318_/X _1323_/C _1327_/Y _1328_/Y _1331_/X VGND VGND VPWR VPWR _2144_/D
+ sky130_fd_sc_hd__a41oi_4
X_1567_ _1569_/A _2189_/Q _1562_/C VGND VGND VPWR VPWR _1568_/D sky130_fd_sc_hd__a21o_4
XFILLER_58_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1636_ _1619_/Y _1621_/B _1293_/X VGND VGND VPWR VPWR _1636_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_58_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2119_ _2025_/CLK _1824_/Y VGND VGND VPWR VPWR _1821_/B sky130_fd_sc_hd__dfxtp_4
X_1498_ _1426_/A _1486_/Y _2146_/Q _1493_/X VGND VGND VPWR VPWR _1498_/Y sky130_fd_sc_hd__nand4_4
XFILLER_22_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_15_0_addressalyzerBlock.SPI_CLK clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2052_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1421_ _1421_/A VGND VGND VPWR VPWR _1421_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1283_ _1291_/A VGND VGND VPWR VPWR _1306_/A sky130_fd_sc_hd__buf_2
XFILLER_36_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1352_ _1164_/X _2040_/D _1172_/X VGND VGND VPWR VPWR _1352_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_63_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0998_ _2247_/Q _0998_/B VGND VGND VPWR VPWR _0998_/X sky130_fd_sc_hd__or2_4
X_1619_ _1607_/X _1646_/C VGND VGND VPWR VPWR _1619_/Y sky130_fd_sc_hd__nor2_4
XFILLER_27_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1970_ _1971_/A _1960_/X _1969_/Y VGND VGND VPWR VPWR _1970_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1335_ _1291_/X _1219_/B _1330_/X VGND VGND VPWR VPWR _1335_/X sky130_fd_sc_hd__a21o_4
X_1404_ _2070_/Q VGND VGND VPWR VPWR _1404_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1197_ _1197_/A VGND VGND VPWR VPWR _1362_/A sky130_fd_sc_hd__buf_2
X_1266_ _1264_/Y _1188_/X _1265_/Y VGND VGND VPWR VPWR _1266_/Y sky130_fd_sc_hd__a21oi_4
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1051_ _1178_/A VGND VGND VPWR VPWR _1052_/B sky130_fd_sc_hd__buf_2
XFILLER_38_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1120_ _1109_/A VGND VGND VPWR VPWR _1120_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1884_ _1765_/Y _1867_/A _1883_/Y VGND VGND VPWR VPWR _2093_/D sky130_fd_sc_hd__o21ai_4
XFILLER_18_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1953_ _1356_/Y _1949_/X _1316_/A _1950_/X VGND VGND VPWR VPWR _1953_/X sky130_fd_sc_hd__a2bb2o_4
X_1318_ _1282_/B VGND VGND VPWR VPWR _1318_/X sky130_fd_sc_hd__buf_2
XFILLER_64_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1249_ _1248_/Y _1209_/A _1272_/B VGND VGND VPWR VPWR _1249_/X sky130_fd_sc_hd__a21o_4
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2221_ _2231_/CLK _1375_/Y VGND VGND VPWR VPWR _1374_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2152_ _2218_/CLK _2152_/D VGND VGND VPWR VPWR _2152_/Q sky130_fd_sc_hd__dfxtp_4
X_1034_ _0996_/X _1004_/X _1034_/C VGND VGND VPWR VPWR _1034_/Y sky130_fd_sc_hd__nand3_4
X_1103_ _2236_/Q VGND VGND VPWR VPWR _1109_/A sky130_fd_sc_hd__buf_2
X_2083_ _2085_/CLK _2083_/D VGND VGND VPWR VPWR _2083_/Q sky130_fd_sc_hd__dfxtp_4
X_1867_ _1867_/A _1767_/B _1867_/C VGND VGND VPWR VPWR _1867_/Y sky130_fd_sc_hd__nand3_4
X_1936_ _1112_/Y _1934_/Y _1733_/D _1462_/Y _1935_/Y VGND VGND VPWR VPWR _1936_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1798_ _1797_/Y _1807_/A _1376_/A _1791_/Y _2131_/Q VGND VGND VPWR VPWR _1798_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_44_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1721_ _1767_/C _1412_/A _1161_/A _1720_/Y VGND VGND VPWR VPWR _1721_/X sky130_fd_sc_hd__a211o_4
X_1652_ _1648_/X _1649_/A _1649_/C _1649_/D _1040_/A VGND VGND VPWR VPWR _1652_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1583_ _1583_/A _1583_/B _2173_/Q _2174_/Q VGND VGND VPWR VPWR _1583_/Y sky130_fd_sc_hd__nand4_4
X_2204_ _2211_/CLK _2204_/D VGND VGND VPWR VPWR _2204_/Q sky130_fd_sc_hd__dfxtp_4
X_2135_ _2137_/CLK _1761_/Y VGND VGND VPWR VPWR _1760_/C sky130_fd_sc_hd__dfxtp_4
X_1017_ _1020_/A _0996_/X _1016_/X VGND VGND VPWR VPWR _1017_/Y sky130_fd_sc_hd__o21ai_4
X_2066_ _2228_/CLK _2066_/D VGND VGND VPWR VPWR _1490_/A sky130_fd_sc_hd__dfxtp_4
X_1919_ _1112_/Y _1916_/X _1918_/Y VGND VGND VPWR VPWR _2081_/D sky130_fd_sc_hd__o21ai_4
XFILLER_57_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1704_ _1704_/A ID_fromClient VGND VGND VPWR VPWR _2145_/D sky130_fd_sc_hd__and2_4
X_1566_ _1564_/X SPI_CLK_RESET_N _1570_/A VGND VGND VPWR VPWR _2191_/D sky130_fd_sc_hd__and3_4
X_1635_ _1584_/C _1632_/Y _1634_/Y VGND VGND VPWR VPWR _1635_/Y sky130_fd_sc_hd__a21oi_4
X_1497_ _1495_/Y _1496_/Y _1446_/X VGND VGND VPWR VPWR _2213_/D sky130_fd_sc_hd__a21oi_4
X_2118_ _2025_/CLK _2118_/D VGND VGND VPWR VPWR _1826_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_39_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2049_ _2211_/CLK _2049_/D VGND VGND VPWR VPWR _2049_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_13_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1420_ _1420_/A _1397_/B _1420_/C VGND VGND VPWR VPWR _1420_/Y sky130_fd_sc_hd__nand3_4
X_1351_ _2088_/Q VGND VGND VPWR VPWR _1351_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1282_ _1282_/A _1282_/B _1282_/C VGND VGND VPWR VPWR _1291_/A sky130_fd_sc_hd__nand3_4
XFILLER_59_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1618_ _1583_/Y VGND VGND VPWR VPWR _1646_/C sky130_fd_sc_hd__buf_2
X_0997_ _0995_/A VGND VGND VPWR VPWR _0998_/B sky130_fd_sc_hd__buf_2
X_1549_ _1549_/A VGND VGND VPWR VPWR _1549_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_1_0_addressalyzerBlock.SPI_CLK clkbuf_3_1_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_4_3_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_24_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1403_ _1402_/Y _1189_/A _1190_/X _1153_/A _1366_/A VGND VGND VPWR VPWR _1403_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1265_ _1790_/A _1243_/B _1243_/C VGND VGND VPWR VPWR _1265_/Y sky130_fd_sc_hd__nor3_4
X_1334_ _1217_/X _1344_/A _1298_/C VGND VGND VPWR VPWR _1334_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_51_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1196_ _1311_/A VGND VGND VPWR VPWR _1196_/X sky130_fd_sc_hd__buf_2
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_0_0_m1_clk_local clkbuf_2_1_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_3_1_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1050_ _1086_/A _1049_/X VGND VGND VPWR VPWR _1052_/A sky130_fd_sc_hd__nor2_4
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1883_ _1864_/Y _1899_/B _2037_/D VGND VGND VPWR VPWR _1883_/Y sky130_fd_sc_hd__nand3_4
XFILLER_14_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1952_ _1487_/Y _1949_/X _1112_/A _1950_/X VGND VGND VPWR VPWR _2065_/D sky130_fd_sc_hd__a2bb2o_4
X_1248_ _1834_/C VGND VGND VPWR VPWR _1248_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1317_ _1215_/A _1071_/X _1313_/Y _1316_/Y _1278_/Y VGND VGND VPWR VPWR _1317_/Y
+ sky130_fd_sc_hd__o32ai_4
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1179_ _1178_/Y VGND VGND VPWR VPWR _1179_/X sky130_fd_sc_hd__buf_2
XFILLER_24_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1102_ _1102_/A VGND VGND VPWR VPWR _1678_/A sky130_fd_sc_hd__buf_2
X_2220_ _2231_/CLK _2220_/D VGND VGND VPWR VPWR _1400_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2151_ _2218_/CLK _1698_/X VGND VGND VPWR VPWR _2151_/Q sky130_fd_sc_hd__dfxtp_4
X_2082_ _2085_/CLK _2082_/D VGND VGND VPWR VPWR ID_toHost sky130_fd_sc_hd__dfxtp_4
XFILLER_61_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1033_ _1029_/Y _1030_/X _1032_/Y VGND VGND VPWR VPWR _1033_/Y sky130_fd_sc_hd__a21oi_4
X_1797_ _1402_/Y _1803_/A _1787_/Y VGND VGND VPWR VPWR _1797_/Y sky130_fd_sc_hd__nor3_4
X_1866_ _1864_/Y VGND VGND VPWR VPWR _1867_/A sky130_fd_sc_hd__buf_2
X_1935_ _1927_/Y _1504_/X VGND VGND VPWR VPWR _1935_/Y sky130_fd_sc_hd__nand2_4
XFILLER_21_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1651_ _2173_/Q _1649_/X _1650_/Y VGND VGND VPWR VPWR _1651_/X sky130_fd_sc_hd__o21a_4
X_1720_ _1154_/X _1719_/Y VGND VGND VPWR VPWR _1720_/Y sky130_fd_sc_hd__nor2_4
X_1582_ _1578_/Y _1579_/Y _1642_/B _1581_/Y VGND VGND VPWR VPWR _1583_/B sky130_fd_sc_hd__nor4_4
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2203_ _2211_/CLK _1528_/X VGND VGND VPWR VPWR _2203_/Q sky130_fd_sc_hd__dfxtp_4
X_2134_ _2137_/CLK _2134_/D VGND VGND VPWR VPWR _1763_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_19_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2065_ _2224_/CLK _2065_/D VGND VGND VPWR VPWR _2065_/Q sky130_fd_sc_hd__dfxtp_4
X_1016_ _2245_/Q _1020_/B VGND VGND VPWR VPWR _1016_/X sky130_fd_sc_hd__or2_4
XFILLER_34_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1849_ _1212_/Y _1779_/B VGND VGND VPWR VPWR _1850_/A sky130_fd_sc_hd__xor2_4
XFILLER_1_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1918_ _1916_/X _1917_/X _2081_/Q VGND VGND VPWR VPWR _1918_/Y sky130_fd_sc_hd__nand3_4
XFILLER_57_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1634_ _1607_/X _1584_/B _1584_/C _1646_/C _1958_/A VGND VGND VPWR VPWR _1634_/Y
+ sky130_fd_sc_hd__o41ai_4
X_1703_ _1704_/A _1703_/B VGND VGND VPWR VPWR _2146_/D sky130_fd_sc_hd__and2_4
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1565_ _1565_/A VGND VGND VPWR VPWR _1570_/A sky130_fd_sc_hd__inv_2
X_1496_ _1426_/Y _2213_/Q VGND VGND VPWR VPWR _1496_/Y sky130_fd_sc_hd__nand2_4
X_2117_ _2025_/CLK _2117_/D VGND VGND VPWR VPWR _1726_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_54_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2048_ _2211_/CLK _2056_/Q VGND VGND VPWR VPWR _2048_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1281_ _1280_/Y VGND VGND VPWR VPWR _1282_/C sky130_fd_sc_hd__inv_2
X_1350_ HASH_LED _1154_/X _1166_/X _1349_/Y VGND VGND VPWR VPWR _1350_/X sky130_fd_sc_hd__a211o_4
XFILLER_36_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0996_ _0996_/A VGND VGND VPWR VPWR _0996_/X sky130_fd_sc_hd__buf_2
X_1617_ _1616_/X _1675_/B _1604_/A VGND VGND VPWR VPWR _2181_/D sky130_fd_sc_hd__and3_4
XFILLER_54_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1479_ _1474_/X _1476_/Y _1478_/Y VGND VGND VPWR VPWR _1479_/X sky130_fd_sc_hd__a21o_4
XFILLER_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1548_ _0995_/A _1455_/D VGND VGND VPWR VPWR _1549_/A sky130_fd_sc_hd__nand2_4
XFILLER_50_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1402_ _1810_/A VGND VGND VPWR VPWR _1402_/Y sky130_fd_sc_hd__inv_2
X_1264_ _1088_/X _1262_/Y _1263_/X VGND VGND VPWR VPWR _1264_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1333_ _1969_/D _1123_/X _1133_/X VGND VGND VPWR VPWR _1333_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_51_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1195_ _1201_/B VGND VGND VPWR VPWR _1195_/X sky130_fd_sc_hd__buf_2
XFILLER_32_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1882_ _1762_/Y _1867_/A _1881_/Y VGND VGND VPWR VPWR _2094_/D sky130_fd_sc_hd__o21ai_4
XFILLER_14_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1951_ _1490_/Y _1949_/X _1894_/A _1950_/X VGND VGND VPWR VPWR _2066_/D sky130_fd_sc_hd__a2bb2o_4
X_1247_ _1203_/Y _2115_/Q _1209_/X VGND VGND VPWR VPWR _1247_/Y sky130_fd_sc_hd__a21oi_4
X_1178_ _1178_/A VGND VGND VPWR VPWR _1178_/Y sky130_fd_sc_hd__inv_2
X_1316_ _1316_/A VGND VGND VPWR VPWR _1316_/Y sky130_fd_sc_hd__inv_2
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1032_ _2219_/Q _1003_/A _1031_/X VGND VGND VPWR VPWR _1032_/Y sky130_fd_sc_hd__o21ai_4
X_1101_ _1098_/A VGND VGND VPWR VPWR _1102_/A sky130_fd_sc_hd__buf_2
X_2150_ _2194_/CLK _1699_/X VGND VGND VPWR VPWR _2150_/Q sky130_fd_sc_hd__dfxtp_4
X_2081_ _2213_/CLK _2081_/D VGND VGND VPWR VPWR _2081_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_61_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1934_ _1896_/Y VGND VGND VPWR VPWR _1934_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1796_ _1796_/A _1796_/B VGND VGND VPWR VPWR _1796_/Y sky130_fd_sc_hd__nor2_4
X_1865_ _1864_/Y VGND VGND VPWR VPWR _1865_/X sky130_fd_sc_hd__buf_2
XFILLER_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1581_ _1668_/A _1581_/B _2166_/Q _2167_/Q VGND VGND VPWR VPWR _1581_/Y sky130_fd_sc_hd__nand4_4
X_1650_ _1649_/C _1642_/Y _1649_/D _2173_/Q _1040_/A VGND VGND VPWR VPWR _1650_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_11_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2202_ _2211_/CLK _1530_/X VGND VGND VPWR VPWR _2202_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1015_ _1013_/Y _1003_/X _1014_/Y VGND VGND VPWR VPWR _2246_/D sky130_fd_sc_hd__a21oi_4
X_2064_ _2224_/CLK _1953_/X VGND VGND VPWR VPWR _2064_/Q sky130_fd_sc_hd__dfxtp_4
X_2133_ _2137_/CLK _2133_/D VGND VGND VPWR VPWR _1767_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_19_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1917_ _1917_/A VGND VGND VPWR VPWR _1917_/X sky130_fd_sc_hd__buf_2
X_1848_ _1847_/X VGND VGND VPWR VPWR _1848_/Y sky130_fd_sc_hd__inv_2
X_1779_ _1779_/A _1779_/B _1776_/Y _1832_/C VGND VGND VPWR VPWR _1840_/B sky130_fd_sc_hd__nand4_4
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_1_0_addressalyzerBlock.SPI_CLK clkbuf_4_1_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2085_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_16_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1564_ _1562_/Y _1563_/A _1563_/Y VGND VGND VPWR VPWR _1564_/X sky130_fd_sc_hd__a21o_4
X_1633_ _1633_/A VGND VGND VPWR VPWR _1958_/A sky130_fd_sc_hd__buf_2
X_1702_ _1701_/A _1702_/B VGND VGND VPWR VPWR _1702_/Y sky130_fd_sc_hd__nand2_4
XFILLER_39_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1495_ _1495_/A _1426_/A _2146_/Q VGND VGND VPWR VPWR _1495_/Y sky130_fd_sc_hd__nand3_4
X_2116_ _2115_/CLK _1833_/Y VGND VGND VPWR VPWR _2116_/Q sky130_fd_sc_hd__dfxtp_4
X_2047_ _2058_/CLK _2047_/D VGND VGND VPWR VPWR _2047_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_54_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_6_0_addressalyzerBlock.SPI_CLK clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
X_1280_ _1280_/A _1064_/Y VGND VGND VPWR VPWR _1280_/Y sky130_fd_sc_hd__nor2_4
XFILLER_48_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0995_ _0995_/A VGND VGND VPWR VPWR _0996_/A sky130_fd_sc_hd__inv_2
XFILLER_59_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1616_ _1608_/Y _1621_/C _1587_/A _1587_/D _2181_/Q VGND VGND VPWR VPWR _1616_/X
+ sky130_fd_sc_hd__a41o_4
X_1547_ _1544_/Y _1545_/Y _1546_/Y VGND VGND VPWR VPWR _2195_/D sky130_fd_sc_hd__a21oi_4
X_1478_ _1477_/Y _1397_/B _1223_/B VGND VGND VPWR VPWR _1478_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_35_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1401_ _1343_/X _1399_/Y _1400_/Y VGND VGND VPWR VPWR _2220_/D sky130_fd_sc_hd__o21ai_4
X_1263_ _1263_/A _1178_/Y VGND VGND VPWR VPWR _1263_/X sky130_fd_sc_hd__or2_4
X_1194_ _1048_/D VGND VGND VPWR VPWR _1201_/B sky130_fd_sc_hd__buf_2
X_1332_ _1318_/X _1323_/C _1327_/Y _1328_/Y _1331_/X VGND VGND VPWR VPWR _2224_/D
+ sky130_fd_sc_hd__a41oi_4
XFILLER_51_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1950_ _1943_/A VGND VGND VPWR VPWR _1950_/X sky130_fd_sc_hd__buf_2
X_1881_ _1871_/X _1899_/B _2038_/D VGND VGND VPWR VPWR _1881_/Y sky130_fd_sc_hd__nand3_4
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1315_ _1314_/X _1306_/A _1215_/A VGND VGND VPWR VPWR _1315_/Y sky130_fd_sc_hd__o21ai_4
X_1246_ _1153_/Y _1244_/Y _1245_/X VGND VGND VPWR VPWR _1246_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_2_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1177_ _1156_/Y _1162_/Y _1176_/Y VGND VGND VPWR VPWR _1177_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_24_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1031_ _1008_/A VGND VGND VPWR VPWR _1031_/X sky130_fd_sc_hd__buf_2
XFILLER_34_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1100_ _1094_/Y _1096_/Y _1099_/X VGND VGND VPWR VPWR _2238_/D sky130_fd_sc_hd__a21oi_4
X_2080_ _2213_/CLK _2080_/D VGND VGND VPWR VPWR HASH_LED sky130_fd_sc_hd__dfxtp_4
X_1933_ _1927_/Y _1341_/C _2074_/Q _1185_/A _1932_/Y VGND VGND VPWR VPWR _2074_/D
+ sky130_fd_sc_hd__a32o_4
X_1795_ _1795_/A _1799_/B VGND VGND VPWR VPWR _1796_/B sky130_fd_sc_hd__nor2_4
X_1864_ _1864_/A VGND VGND VPWR VPWR _1864_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1229_ _1229_/A _1229_/B VGND VGND VPWR VPWR _2232_/D sky130_fd_sc_hd__nand2_4
XFILLER_12_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1580_ _2168_/Q _1580_/B VGND VGND VPWR VPWR _1642_/B sky130_fd_sc_hd__nand2_4
XFILLER_7_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2132_ _2124_/CLK _1796_/Y VGND VGND VPWR VPWR _1192_/A sky130_fd_sc_hd__dfxtp_4
X_2201_ _2211_/CLK _2201_/D VGND VGND VPWR VPWR _2201_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1014_ _2230_/Q _1004_/X _1008_/X VGND VGND VPWR VPWR _1014_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2063_ _2224_/CLK _1954_/X VGND VGND VPWR VPWR _1388_/A sky130_fd_sc_hd__dfxtp_4
X_1847_ _1847_/A _1847_/B VGND VGND VPWR VPWR _1847_/X sky130_fd_sc_hd__xor2_4
X_1916_ _1915_/Y VGND VGND VPWR VPWR _1916_/X sky130_fd_sc_hd__buf_2
X_1778_ _1777_/Y VGND VGND VPWR VPWR _1832_/C sky130_fd_sc_hd__inv_2
XFILLER_17_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1701_ _1701_/A _1688_/Y VGND VGND VPWR VPWR _1701_/Y sky130_fd_sc_hd__nand2_4
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1563_ _1563_/A _1570_/C VGND VGND VPWR VPWR _1563_/Y sky130_fd_sc_hd__nor2_4
X_1632_ _1608_/Y VGND VGND VPWR VPWR _1632_/Y sky130_fd_sc_hd__inv_2
X_1494_ _1486_/Y _1493_/X _1061_/D VGND VGND VPWR VPWR _1495_/A sky130_fd_sc_hd__a21o_4
XFILLER_3_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2115_ _2115_/CLK _1837_/Y VGND VGND VPWR VPWR _2115_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2046_ _2044_/CLK _2046_/D VGND VGND VPWR VPWR _2046_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_5_0_m1_clk_local clkbuf_3_4_0_m1_clk_local/A VGND VGND VPWR VPWR _2029_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1477_ _2105_/Q VGND VGND VPWR VPWR _1477_/Y sky130_fd_sc_hd__inv_2
X_1615_ _1609_/B VGND VGND VPWR VPWR _1621_/C sky130_fd_sc_hd__buf_2
XFILLER_5_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1546_ _1455_/Y _1456_/Y VGND VGND VPWR VPWR _1546_/Y sky130_fd_sc_hd__nand2_4
XFILLER_54_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2029_ _2029_/CLK _2029_/D VGND VGND VPWR VPWR MACRO_RD_SELECT sky130_fd_sc_hd__dfxtp_4
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1400_ _1274_/A _1400_/B VGND VGND VPWR VPWR _1400_/Y sky130_fd_sc_hd__nand2_4
X_1331_ _1291_/X _1329_/X _1330_/X VGND VGND VPWR VPWR _1331_/X sky130_fd_sc_hd__a21o_4
XFILLER_5_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1193_ _1181_/Y _1188_/X _1192_/Y VGND VGND VPWR VPWR _1193_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1262_ _1253_/Y _1254_/Y _1261_/Y VGND VGND VPWR VPWR _1262_/Y sky130_fd_sc_hd__a21oi_4
X_1529_ _2202_/Q _1526_/X _1521_/X VGND VGND VPWR VPWR _1529_/X sky130_fd_sc_hd__o21a_4
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1880_ _1759_/Y _1867_/A _1879_/Y VGND VGND VPWR VPWR _1880_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_14_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1314_ _1308_/X _1451_/A _1313_/Y VGND VGND VPWR VPWR _1314_/X sky130_fd_sc_hd__o21a_4
X_1245_ _1195_/X _1813_/A _1196_/X _1473_/C VGND VGND VPWR VPWR _1245_/X sky130_fd_sc_hd__a211o_4
XFILLER_2_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1176_ _1168_/Y _1174_/Y _1175_/X VGND VGND VPWR VPWR _1176_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_24_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1030_ _1004_/A VGND VGND VPWR VPWR _1030_/X sky130_fd_sc_hd__buf_2
XFILLER_61_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1932_ _1748_/Y VGND VGND VPWR VPWR _1932_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1863_ _1396_/C _1005_/Y _1152_/D _2217_/Q VGND VGND VPWR VPWR _1864_/A sky130_fd_sc_hd__and4_4
X_1794_ _2131_/Q _1807_/B _1807_/A _1791_/Y VGND VGND VPWR VPWR _1799_/B sky130_fd_sc_hd__nand4_4
XFILLER_6_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1228_ _1274_/A _1228_/B VGND VGND VPWR VPWR _1229_/B sky130_fd_sc_hd__nand2_4
XFILLER_52_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1159_ _1170_/A VGND VGND VPWR VPWR _1159_/X sky130_fd_sc_hd__buf_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2131_ _2124_/CLK _2131_/D VGND VGND VPWR VPWR _2131_/Q sky130_fd_sc_hd__dfxtp_4
X_2200_ _2194_/CLK _2200_/D VGND VGND VPWR VPWR _2200_/Q sky130_fd_sc_hd__dfxtp_4
X_2062_ _2224_/CLK _1955_/X VGND VGND VPWR VPWR _1482_/A sky130_fd_sc_hd__dfxtp_4
X_1013_ _2245_/Q _0996_/X _1012_/X VGND VGND VPWR VPWR _1013_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_4_6_0_addressalyzerBlock.SPI_CLK clkbuf_4_7_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2228_/CLK sky130_fd_sc_hd__clkbuf_1
X_1846_ _1846_/A _1845_/Y VGND VGND VPWR VPWR _1846_/Y sky130_fd_sc_hd__xnor2_4
X_1777_ _1777_/A _1843_/A VGND VGND VPWR VPWR _1777_/Y sky130_fd_sc_hd__nand2_4
X_1915_ _1914_/Y VGND VGND VPWR VPWR _1915_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1631_ _1624_/D _1584_/Y _1630_/Y VGND VGND VPWR VPWR _2178_/D sky130_fd_sc_hd__o21a_4
X_1700_ _1704_/A MOSI_fromHost VGND VGND VPWR VPWR _1700_/X sky130_fd_sc_hd__and2_4
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1562_ _1569_/A _2189_/Q _1562_/C VGND VGND VPWR VPWR _1562_/Y sky130_fd_sc_hd__nand3_4
X_1493_ _1488_/X _1489_/Y _1491_/Y _1492_/Y VGND VGND VPWR VPWR _1493_/X sky130_fd_sc_hd__and4_4
X_2114_ _2115_/CLK _1839_/X VGND VGND VPWR VPWR _1770_/A sky130_fd_sc_hd__dfxtp_4
X_2045_ _2044_/CLK _2053_/Q VGND VGND VPWR VPWR _2045_/Q sky130_fd_sc_hd__dfxtp_4
X_1829_ _1834_/A _1834_/B _1834_/C _1776_/Y VGND VGND VPWR VPWR _1829_/X sky130_fd_sc_hd__and4_4
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1614_ _1595_/A _1604_/A _1613_/Y VGND VGND VPWR VPWR _1614_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1476_ _1203_/Y _1840_/A _1209_/A VGND VGND VPWR VPWR _1476_/Y sky130_fd_sc_hd__a21oi_4
X_1545_ _0998_/B _1455_/C _1455_/D VGND VGND VPWR VPWR _1545_/Y sky130_fd_sc_hd__nand3_4
XFILLER_54_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2028_ _2189_/CLK _2028_/D VGND VGND VPWR VPWR DATA_TO_HASH[7] sky130_fd_sc_hd__dfxtp_4
XFILLER_42_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1330_ _1330_/A VGND VGND VPWR VPWR _1330_/X sky130_fd_sc_hd__buf_2
X_1261_ _1257_/Y _1260_/Y _1175_/X VGND VGND VPWR VPWR _1261_/Y sky130_fd_sc_hd__a21oi_4
X_1192_ _1192_/A _1243_/B _1243_/C VGND VGND VPWR VPWR _1192_/Y sky130_fd_sc_hd__nor3_4
XFILLER_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1528_ _2202_/Q _1525_/X _1527_/X VGND VGND VPWR VPWR _1528_/X sky130_fd_sc_hd__o21a_4
XFILLER_19_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1459_ _1159_/X _2065_/Q _1161_/A VGND VGND VPWR VPWR _1459_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1244_ _1242_/Y _1188_/X _1243_/Y VGND VGND VPWR VPWR _1244_/Y sky130_fd_sc_hd__a21oi_4
X_1313_ _1310_/X _1313_/B _1312_/X VGND VGND VPWR VPWR _1313_/Y sky130_fd_sc_hd__nand3_4
XFILLER_2_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1175_ _2144_/Q VGND VGND VPWR VPWR _1175_/X sky130_fd_sc_hd__buf_2
XFILLER_55_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1793_ _1192_/A VGND VGND VPWR VPWR _1795_/A sky130_fd_sc_hd__inv_2
X_1862_ _1857_/A _2101_/Q VGND VGND VPWR VPWR _1862_/X sky130_fd_sc_hd__xor2_4
X_1931_ _1927_/Y _1341_/C _2075_/Q _1185_/A _1930_/Y VGND VGND VPWR VPWR _2075_/D
+ sky130_fd_sc_hd__a32o_4
X_1227_ _1480_/A VGND VGND VPWR VPWR _1274_/A sky130_fd_sc_hd__buf_2
XFILLER_25_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1158_ _1171_/A VGND VGND VPWR VPWR _1170_/A sky130_fd_sc_hd__buf_2
XFILLER_40_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1089_ _1088_/X VGND VGND VPWR VPWR _1089_/X sky130_fd_sc_hd__buf_2
XFILLER_12_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_11_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2218_/CLK sky130_fd_sc_hd__clkbuf_1
X_2130_ _2124_/CLK _2130_/D VGND VGND VPWR VPWR _1790_/A sky130_fd_sc_hd__dfxtp_4
X_1012_ _2246_/Q _1020_/B VGND VGND VPWR VPWR _1012_/X sky130_fd_sc_hd__or2_4
XFILLER_19_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2061_ _2228_/CLK _1956_/X VGND VGND VPWR VPWR _1483_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_34_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1914_ _1038_/A _1310_/A _1886_/C _1909_/X VGND VGND VPWR VPWR _1914_/Y sky130_fd_sc_hd__nor4_4
XFILLER_22_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1776_ _1775_/Y VGND VGND VPWR VPWR _1776_/Y sky130_fd_sc_hd__inv_2
X_1845_ _2109_/Q _1834_/A _1834_/B _1834_/C VGND VGND VPWR VPWR _1845_/Y sky130_fd_sc_hd__nand4_4
XFILLER_8_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1630_ _1621_/B _1619_/Y _1621_/C _1624_/D _1040_/A VGND VGND VPWR VPWR _1630_/Y
+ sky130_fd_sc_hd__a41oi_4
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1561_ _1560_/X VGND VGND VPWR VPWR _2192_/D sky130_fd_sc_hd__inv_2
X_1492_ _1126_/B _1482_/A _2235_/Q _1389_/B VGND VGND VPWR VPWR _1492_/Y sky130_fd_sc_hd__a22oi_4
X_2044_ _2044_/CLK DATA_AVAILABLE VGND VGND VPWR VPWR _2044_/Q sky130_fd_sc_hd__dfxtp_4
X_2113_ _2025_/CLK _2113_/D VGND VGND VPWR VPWR _1475_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_30_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1828_ _1371_/X _1774_/C _1774_/D VGND VGND VPWR VPWR _1834_/A sky130_fd_sc_hd__nor3_4
X_1759_ _1504_/X _1445_/A _1902_/A VGND VGND VPWR VPWR _1759_/Y sky130_fd_sc_hd__nand3_4
XFILLER_54_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1613_ _1595_/A _1604_/A _1031_/X VGND VGND VPWR VPWR _1613_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1544_ _1544_/A VGND VGND VPWR VPWR _1544_/Y sky130_fd_sc_hd__inv_2
X_1475_ _1475_/A VGND VGND VPWR VPWR _1840_/A sky130_fd_sc_hd__inv_2
XFILLER_39_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2027_ _2029_/CLK _2027_/D VGND VGND VPWR VPWR DATA_TO_HASH[6] sky130_fd_sc_hd__dfxtp_4
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1191_ _1190_/X VGND VGND VPWR VPWR _1243_/C sky130_fd_sc_hd__buf_2
X_1260_ _1258_/Y _1170_/X _1259_/Y VGND VGND VPWR VPWR _1260_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_36_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_1_0_m1_clk_local clkbuf_3_1_0_m1_clk_local/A VGND VGND VPWR VPWR _2171_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_1527_ _2203_/Q _1526_/X _1521_/X VGND VGND VPWR VPWR _1527_/X sky130_fd_sc_hd__o21a_4
X_1458_ _1455_/Y _1458_/B VGND VGND VPWR VPWR _2215_/D sky130_fd_sc_hd__nor2_4
X_1389_ _1412_/A _1389_/B VGND VGND VPWR VPWR _1389_/Y sky130_fd_sc_hd__nor2_4
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1243_ _2131_/Q _1243_/B _1243_/C VGND VGND VPWR VPWR _1243_/Y sky130_fd_sc_hd__nor3_4
X_1312_ _1201_/B VGND VGND VPWR VPWR _1312_/X sky130_fd_sc_hd__buf_2
XFILLER_37_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1174_ _1169_/Y _1170_/X _1173_/Y VGND VGND VPWR VPWR _1174_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_32_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1930_ _1930_/A VGND VGND VPWR VPWR _1930_/Y sky130_fd_sc_hd__inv_2
X_1792_ _2131_/Q _1807_/B _1807_/A _1791_/Y _1192_/A VGND VGND VPWR VPWR _1796_/A
+ sky130_fd_sc_hd__a41oi_4
X_1861_ _2102_/Q _1860_/Y VGND VGND VPWR VPWR _1861_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_6_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1226_ _1226_/A VGND VGND VPWR VPWR _1480_/A sky130_fd_sc_hd__buf_2
X_1157_ _2142_/Q VGND VGND VPWR VPWR _1171_/A sky130_fd_sc_hd__inv_2
X_1088_ _1052_/B VGND VGND VPWR VPWR _1088_/X sky130_fd_sc_hd__buf_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2060_ _2052_/CLK DATA_FROM_HASH[7] VGND VGND VPWR VPWR _2052_/D sky130_fd_sc_hd__dfxtp_4
X_1011_ _0995_/A VGND VGND VPWR VPWR _1020_/B sky130_fd_sc_hd__buf_2
XFILLER_8_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1913_ _1894_/Y _1909_/X _1905_/X _1255_/Y _1910_/X VGND VGND VPWR VPWR _2082_/D
+ sky130_fd_sc_hd__o32ai_4
X_1775_ _1846_/A _2109_/Q VGND VGND VPWR VPWR _1775_/Y sky130_fd_sc_hd__nand2_4
X_1844_ _1844_/A VGND VGND VPWR VPWR _2111_/D sky130_fd_sc_hd__inv_2
XFILLER_8_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2189_ _2189_/CLK _2189_/D VGND VGND VPWR VPWR _2189_/Q sky130_fd_sc_hd__dfxtp_4
X_1209_ _1209_/A VGND VGND VPWR VPWR _1209_/X sky130_fd_sc_hd__buf_2
XFILLER_25_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1560_ _2192_/Q _1565_/A _1559_/Y VGND VGND VPWR VPWR _1560_/X sky130_fd_sc_hd__a21o_4
XFILLER_33_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2112_ _2025_/CLK _2112_/D VGND VGND VPWR VPWR _1777_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_39_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1491_ _1120_/Y _2064_/Q _1076_/B _1490_/Y VGND VGND VPWR VPWR _1491_/Y sky130_fd_sc_hd__a22oi_4
X_2043_ _2058_/CLK _2044_/Q VGND VGND VPWR VPWR _2043_/Q sky130_fd_sc_hd__dfxtp_4
X_1827_ _1825_/B _1827_/B VGND VGND VPWR VPWR _2117_/D sky130_fd_sc_hd__xor2_4
X_1758_ _1739_/X _1756_/Y _1757_/Y VGND VGND VPWR VPWR _2136_/D sky130_fd_sc_hd__o21ai_4
X_1689_ _1704_/A _1688_/Y _2148_/Q VGND VGND VPWR VPWR _1689_/X sky130_fd_sc_hd__and3_4
XFILLER_57_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_2_0_addressalyzerBlock.SPI_CLK clkbuf_2_3_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_53_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1474_ _1470_/Y _1471_/X _1203_/Y _1473_/Y VGND VGND VPWR VPWR _1474_/X sky130_fd_sc_hd__a211o_4
X_1612_ _1611_/Y VGND VGND VPWR VPWR _2183_/D sky130_fd_sc_hd__inv_2
X_1543_ _1524_/Y _2150_/Q _1542_/X VGND VGND VPWR VPWR _1543_/X sky130_fd_sc_hd__o21a_4
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2026_ _2182_/CLK _2026_/D VGND VGND VPWR VPWR DATA_TO_HASH[5] sky130_fd_sc_hd__dfxtp_4
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1190_ _1185_/Y VGND VGND VPWR VPWR _1190_/X sky130_fd_sc_hd__buf_2
XFILLER_39_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1526_ _2156_/Q VGND VGND VPWR VPWR _1526_/X sky130_fd_sc_hd__buf_2
X_1457_ _1456_/Y VGND VGND VPWR VPWR _1458_/B sky130_fd_sc_hd__inv_2
XFILLER_35_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1388_ _1388_/A VGND VGND VPWR VPWR _1389_/B sky130_fd_sc_hd__inv_2
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2009_ _2216_/CLK _1959_/Y VGND VGND VPWR VPWR _1431_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_2_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1311_ _1311_/A VGND VGND VPWR VPWR _1313_/B sky130_fd_sc_hd__buf_2
XFILLER_64_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1242_ _1088_/X _1240_/Y _1241_/X VGND VGND VPWR VPWR _1242_/Y sky130_fd_sc_hd__o21ai_4
X_1173_ _1171_/X _1867_/C _1172_/X VGND VGND VPWR VPWR _1173_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_20_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1509_ _1005_/Y VGND VGND VPWR VPWR _1633_/A sky130_fd_sc_hd__buf_2
XFILLER_55_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1860_ _1857_/A _2101_/Q VGND VGND VPWR VPWR _1860_/Y sky130_fd_sc_hd__nand2_4
XFILLER_52_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1791_ _1791_/A VGND VGND VPWR VPWR _1791_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1225_ _1200_/Y _1210_/Y _1224_/X VGND VGND VPWR VPWR _1229_/A sky130_fd_sc_hd__a21o_4
X_1087_ _1084_/Y _1085_/Y _1086_/X _1049_/X VGND VGND VPWR VPWR _1087_/Y sky130_fd_sc_hd__nor4_4
XFILLER_37_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1156_ _1156_/A _1155_/X VGND VGND VPWR VPWR _1156_/Y sky130_fd_sc_hd__nand2_4
X_1989_ _1228_/B _1003_/A _1969_/A VGND VGND VPWR VPWR _1989_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1010_ _0999_/Y _1003_/X _1009_/Y VGND VGND VPWR VPWR _2247_/D sky130_fd_sc_hd__a21oi_4
XFILLER_34_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1843_ _1843_/A _1832_/B VGND VGND VPWR VPWR _1844_/A sky130_fd_sc_hd__xnor2_4
X_1912_ _1892_/Y _1909_/X _1905_/X _1232_/Y _1910_/X VGND VGND VPWR VPWR _2083_/D
+ sky130_fd_sc_hd__o32ai_4
X_1774_ _1248_/Y _1371_/A _1774_/C _1774_/D VGND VGND VPWR VPWR _1779_/B sky130_fd_sc_hd__nor4_4
X_1208_ _1207_/X VGND VGND VPWR VPWR _1209_/A sky130_fd_sc_hd__buf_2
X_2188_ _2124_/CLK _2188_/D VGND VGND VPWR VPWR _1569_/A sky130_fd_sc_hd__dfxtp_4
X_1139_ _2204_/Q VGND VGND VPWR VPWR _1907_/A sky130_fd_sc_hd__buf_2
XFILLER_0_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1490_ _1490_/A VGND VGND VPWR VPWR _1490_/Y sky130_fd_sc_hd__inv_2
X_2111_ _2115_/CLK _2111_/D VGND VGND VPWR VPWR _1843_/A sky130_fd_sc_hd__dfxtp_4
X_2042_ _2171_/CLK _2098_/Q VGND VGND VPWR VPWR _2036_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_62_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1826_ _1826_/A _1826_/B VGND VGND VPWR VPWR _2118_/D sky130_fd_sc_hd__xor2_4
X_1757_ _1754_/A _1754_/B _1757_/C VGND VGND VPWR VPWR _1757_/Y sky130_fd_sc_hd__nand3_4
X_1688_ _2147_/Q VGND VGND VPWR VPWR _1688_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1611_ _1600_/B _1589_/B _1610_/Y VGND VGND VPWR VPWR _1611_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_8_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1473_ _1820_/A _1473_/B _1473_/C VGND VGND VPWR VPWR _1473_/Y sky130_fd_sc_hd__nor3_4
X_1542_ _2196_/Q _2156_/Q _1535_/X VGND VGND VPWR VPWR _1542_/X sky130_fd_sc_hd__o21a_4
X_2025_ _2025_/CLK _2001_/Q VGND VGND VPWR VPWR DATA_TO_HASH[4] sky130_fd_sc_hd__dfxtp_4
XFILLER_54_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1809_ _1376_/A _1797_/Y VGND VGND VPWR VPWR _2127_/D sky130_fd_sc_hd__xor2_4
XFILLER_49_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1525_ _1524_/Y VGND VGND VPWR VPWR _1525_/X sky130_fd_sc_hd__buf_2
X_1387_ _1355_/A VGND VGND VPWR VPWR _1412_/A sky130_fd_sc_hd__buf_2
X_1456_ _1330_/A _2158_/Q VGND VGND VPWR VPWR _1456_/Y sky130_fd_sc_hd__nor2_4
XFILLER_35_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2008_ _2248_/CLK _2008_/D VGND VGND VPWR VPWR _1449_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1310_ _1310_/A VGND VGND VPWR VPWR _1310_/X sky130_fd_sc_hd__buf_2
X_1241_ _1241_/A _1179_/X VGND VGND VPWR VPWR _1241_/X sky130_fd_sc_hd__or2_4
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1172_ _2143_/Q VGND VGND VPWR VPWR _1172_/X sky130_fd_sc_hd__buf_2
XFILLER_17_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1508_ _1573_/B _2202_/Q _1507_/X VGND VGND VPWR VPWR _1508_/X sky130_fd_sc_hd__o21a_4
X_1439_ _2217_/Q VGND VGND VPWR VPWR _1886_/C sky130_fd_sc_hd__inv_2
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1790_ _1790_/A _2129_/Q VGND VGND VPWR VPWR _1791_/A sky130_fd_sc_hd__nand2_4
X_1224_ _1212_/Y _1209_/X _1272_/B VGND VGND VPWR VPWR _1224_/X sky130_fd_sc_hd__a21o_4
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1086_ _1086_/A VGND VGND VPWR VPWR _1086_/X sky130_fd_sc_hd__buf_2
X_1155_ _1154_/X VGND VGND VPWR VPWR _1155_/X sky130_fd_sc_hd__buf_2
X_1988_ _2247_/Q _0996_/A _1987_/X VGND VGND VPWR VPWR _1988_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_3_0_m1_clk_local clkbuf_2_3_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_3_7_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_2_0_addressalyzerBlock.SPI_CLK clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR clkbuf_4_5_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_19_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1842_ _1777_/A _1841_/Y VGND VGND VPWR VPWR _2112_/D sky130_fd_sc_hd__xnor2_4
X_1773_ _1773_/A _1773_/B _2102_/Q _2101_/Q VGND VGND VPWR VPWR _1774_/D sky130_fd_sc_hd__nand4_4
X_1911_ _1042_/Y _1909_/X _1905_/X _1163_/Y _1910_/X VGND VGND VPWR VPWR _2084_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_6_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1207_ _1344_/B _1207_/B _1344_/C _1344_/D VGND VGND VPWR VPWR _1207_/X sky130_fd_sc_hd__and4_4
X_2187_ _2213_/CLK _1573_/Y VGND VGND VPWR VPWR _1280_/A sky130_fd_sc_hd__dfxtp_4
X_1138_ _1091_/X _1053_/X _1137_/Y VGND VGND VPWR VPWR _1138_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_40_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1069_ _1062_/Y _1069_/B VGND VGND VPWR VPWR _1069_/Y sky130_fd_sc_hd__nand2_4
XFILLER_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2041_ _2025_/CLK _2041_/D VGND VGND VPWR VPWR _2041_/Q sky130_fd_sc_hd__dfxtp_4
X_2110_ _2115_/CLK _1846_/Y VGND VGND VPWR VPWR _1846_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_39_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1825_ _1825_/A _1825_/B VGND VGND VPWR VPWR _1826_/B sky130_fd_sc_hd__and2_4
XFILLER_30_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1756_ _1958_/A _1445_/A _1316_/A VGND VGND VPWR VPWR _1756_/Y sky130_fd_sc_hd__nand3_4
XFILLER_57_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1687_ _1681_/A VGND VGND VPWR VPWR _1704_/A sky130_fd_sc_hd__buf_2
X_2239_ _2051_/CLK _1082_/Y VGND VGND VPWR VPWR _1059_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_21_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1610_ _2181_/Q _1609_/X _1574_/A _1600_/B _1330_/X VGND VGND VPWR VPWR _1610_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1472_ _2121_/Q VGND VGND VPWR VPWR _1820_/A sky130_fd_sc_hd__inv_2
X_1541_ _2196_/Q _1524_/Y _1540_/X VGND VGND VPWR VPWR _1541_/X sky130_fd_sc_hd__o21a_4
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2024_ _2182_/CLK _2024_/D VGND VGND VPWR VPWR DATA_TO_HASH[3] sky130_fd_sc_hd__dfxtp_4
XFILLER_62_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1808_ _1808_/A VGND VGND VPWR VPWR _1808_/Y sky130_fd_sc_hd__inv_2
X_1739_ _1738_/Y VGND VGND VPWR VPWR _1739_/X sky130_fd_sc_hd__buf_2
XFILLER_41_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1524_ _2156_/Q VGND VGND VPWR VPWR _1524_/Y sky130_fd_sc_hd__inv_2
X_1386_ _1382_/X _1385_/Y _2144_/Q VGND VGND VPWR VPWR _1386_/X sky130_fd_sc_hd__a21o_4
X_1455_ _1544_/A _0998_/B _1455_/C _1455_/D VGND VGND VPWR VPWR _1455_/Y sky130_fd_sc_hd__nand4_4
X_2007_ _2218_/CLK _1973_/X VGND VGND VPWR VPWR _1065_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_23_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1240_ _1230_/Y _1231_/Y _1239_/Y VGND VGND VPWR VPWR _1240_/Y sky130_fd_sc_hd__a21oi_4
X_1171_ _1171_/A VGND VGND VPWR VPWR _1171_/X sky130_fd_sc_hd__buf_2
XFILLER_2_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1507_ _1503_/X _1892_/A _1504_/X VGND VGND VPWR VPWR _1507_/X sky130_fd_sc_hd__o21a_4
XFILLER_55_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1369_ _1364_/Y _1397_/B _1369_/C VGND VGND VPWR VPWR _1369_/Y sky130_fd_sc_hd__nand3_4
X_1438_ _1448_/A _1451_/B _1449_/C VGND VGND VPWR VPWR _1438_/Y sky130_fd_sc_hd__nor3_4
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1223_ _1223_/A _1223_/B VGND VGND VPWR VPWR _1272_/B sky130_fd_sc_hd__nand2_4
XFILLER_37_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1154_ _2142_/Q VGND VGND VPWR VPWR _1154_/X sky130_fd_sc_hd__buf_2
XFILLER_52_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1085_ _1149_/A VGND VGND VPWR VPWR _1085_/Y sky130_fd_sc_hd__inv_2
X_1987_ _1987_/A _1020_/B VGND VGND VPWR VPWR _1987_/X sky130_fd_sc_hd__or2_4
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1910_ _1329_/X _1196_/X _1195_/X _1740_/X _1098_/A VGND VGND VPWR VPWR _1910_/X
+ sky130_fd_sc_hd__a41o_4
X_1841_ _1843_/A _1779_/B _1834_/B _1776_/Y VGND VGND VPWR VPWR _1841_/Y sky130_fd_sc_hd__nand4_4
X_1772_ _1772_/A _2105_/Q VGND VGND VPWR VPWR _1774_/C sky130_fd_sc_hd__nand2_4
X_2186_ _2189_/CLK _1598_/Y VGND VGND VPWR VPWR CLK_LED sky130_fd_sc_hd__dfxtp_4
X_1137_ _1091_/X _1105_/A _1089_/X _1125_/D _1957_/C VGND VGND VPWR VPWR _1137_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1206_ _1206_/A VGND VGND VPWR VPWR _1207_/B sky130_fd_sc_hd__inv_2
XFILLER_43_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1068_ _1067_/Y VGND VGND VPWR VPWR _1069_/B sky130_fd_sc_hd__inv_2
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2040_ _2029_/CLK _2040_/D VGND VGND VPWR VPWR _2034_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_62_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1824_ _1821_/B _1824_/B VGND VGND VPWR VPWR _1824_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_30_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1686_ _1697_/A _1987_/A VGND VGND VPWR VPWR _1686_/X sky130_fd_sc_hd__and2_4
X_1755_ _1739_/X _1753_/Y _1754_/Y VGND VGND VPWR VPWR _1755_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_57_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2238_ _2051_/CLK _2238_/D VGND VGND VPWR VPWR _1097_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_53_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2169_ _2171_/CLK _2169_/D VGND VGND VPWR VPWR _1580_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_5_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1540_ _2197_/Q _2156_/Q _1535_/X VGND VGND VPWR VPWR _1540_/X sky130_fd_sc_hd__o21a_4
X_1471_ _2129_/Q _1189_/A _1190_/X _1153_/A _1362_/A VGND VGND VPWR VPWR _1471_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_39_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2023_ _2029_/CLK _1999_/Q VGND VGND VPWR VPWR DATA_TO_HASH[2] sky130_fd_sc_hd__dfxtp_4
X_1807_ _1807_/A _1807_/B VGND VGND VPWR VPWR _1808_/A sky130_fd_sc_hd__xnor2_4
X_1669_ _1581_/B VGND VGND VPWR VPWR _1670_/B sky130_fd_sc_hd__buf_2
X_1738_ _1738_/A VGND VGND VPWR VPWR _1738_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1454_ _1454_/A VGND VGND VPWR VPWR _1454_/Y sky130_fd_sc_hd__inv_2
X_1523_ _1501_/Y _2196_/Q _1522_/X VGND VGND VPWR VPWR _2204_/D sky130_fd_sc_hd__o21a_4
XFILLER_27_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1385_ _1383_/Y _1233_/X _1384_/Y VGND VGND VPWR VPWR _1385_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2006_ _2218_/CLK _2006_/D VGND VGND VPWR VPWR _2006_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_2_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1170_ _1170_/A VGND VGND VPWR VPWR _1170_/X sky130_fd_sc_hd__buf_2
XFILLER_64_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1437_ _1451_/C VGND VGND VPWR VPWR _1449_/C sky130_fd_sc_hd__inv_2
Xclkbuf_4_2_0_addressalyzerBlock.SPI_CLK clkbuf_4_3_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2137_/CLK sky130_fd_sc_hd__clkbuf_1
X_1506_ _1573_/B _2203_/Q _1505_/X VGND VGND VPWR VPWR _2211_/D sky130_fd_sc_hd__o21a_4
X_1368_ _1396_/A _1777_/A _1396_/C VGND VGND VPWR VPWR _1369_/C sky130_fd_sc_hd__nand3_4
X_1299_ _1064_/A _2012_/Q _1894_/A VGND VGND VPWR VPWR _1299_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_23_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_7_0_addressalyzerBlock.SPI_CLK clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1153_ _1153_/A _1197_/A VGND VGND VPWR VPWR _1153_/Y sky130_fd_sc_hd__nor2_4
X_1222_ _1217_/X _1344_/A _1708_/A VGND VGND VPWR VPWR _1223_/B sky130_fd_sc_hd__o21ai_4
X_1084_ _1125_/D VGND VGND VPWR VPWR _1084_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1986_ _2043_/Q _2161_/Q VGND VGND VPWR VPWR IRQ_OUT_toHost sky130_fd_sc_hd__or2_4
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1840_ _1840_/A _1840_/B VGND VGND VPWR VPWR _2113_/D sky130_fd_sc_hd__xor2_4
XFILLER_63_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1771_ _2116_/Q _2115_/Q VGND VGND VPWR VPWR _1780_/B sky130_fd_sc_hd__nand2_4
XFILLER_6_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2185_ _2189_/CLK _2185_/D VGND VGND VPWR VPWR _2185_/Q sky130_fd_sc_hd__dfxtp_4
X_1067_ _1282_/A _1064_/Y _1282_/B VGND VGND VPWR VPWR _1067_/Y sky130_fd_sc_hd__nand3_4
X_1205_ _1047_/A _1048_/D VGND VGND VPWR VPWR _1206_/A sky130_fd_sc_hd__nand2_4
X_1136_ _1132_/Y _1134_/Y _1135_/X VGND VGND VPWR VPWR _1136_/Y sky130_fd_sc_hd__a21oi_4
X_1969_ _1969_/A _2240_/Q _1036_/B _1969_/D VGND VGND VPWR VPWR _1969_/Y sky130_fd_sc_hd__nand4_4
XFILLER_56_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1823_ _1827_/B _1826_/A _1825_/B VGND VGND VPWR VPWR _1824_/B sky130_fd_sc_hd__nand3_4
XFILLER_30_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1685_ _1697_/A IRQ_OUT_fromClient VGND VGND VPWR VPWR _1685_/X sky130_fd_sc_hd__and2_4
X_1754_ _1754_/A _1754_/B _1460_/A VGND VGND VPWR VPWR _1754_/Y sky130_fd_sc_hd__nand3_4
X_2237_ _2228_/CLK _2237_/D VGND VGND VPWR VPWR _1057_/A sky130_fd_sc_hd__dfxtp_4
X_2168_ _2171_/CLK _1667_/Y VGND VGND VPWR VPWR _2168_/Q sky130_fd_sc_hd__dfxtp_4
X_1119_ _1316_/A _1078_/X _1079_/X VGND VGND VPWR VPWR _1119_/Y sky130_fd_sc_hd__a21oi_4
X_2099_ _2091_/CLK _2099_/D VGND VGND VPWR VPWR _1869_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1470_ _1461_/X _1468_/Y _1469_/Y VGND VGND VPWR VPWR _1470_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_5_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2022_ _2189_/CLK _1998_/Q VGND VGND VPWR VPWR DATA_TO_HASH[1] sky130_fd_sc_hd__dfxtp_4
XFILLER_50_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1806_ _1806_/A VGND VGND VPWR VPWR _2129_/D sky130_fd_sc_hd__inv_2
X_1668_ _1668_/A VGND VGND VPWR VPWR _1668_/X sky130_fd_sc_hd__buf_2
X_1599_ _1589_/A VGND VGND VPWR VPWR _1600_/B sky130_fd_sc_hd__buf_2
X_1737_ _1219_/B _1310_/A _1201_/B _2217_/Q VGND VGND VPWR VPWR _1738_/A sky130_fd_sc_hd__and4_4
XFILLER_53_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1453_ _1450_/X _1451_/Y _1452_/Y VGND VGND VPWR VPWR _1454_/A sky130_fd_sc_hd__o21ai_4
XFILLER_4_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1522_ _2215_/Q _1907_/A _1521_/X VGND VGND VPWR VPWR _1522_/X sky130_fd_sc_hd__o21a_4
XFILLER_55_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1384_ _1164_/X _2039_/D _1172_/X VGND VGND VPWR VPWR _1384_/Y sky130_fd_sc_hd__a21oi_4
X_2005_ _2218_/CLK _1976_/Y VGND VGND VPWR VPWR _2006_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_35_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1367_ _1202_/A VGND VGND VPWR VPWR _1396_/C sky130_fd_sc_hd__buf_2
XFILLER_28_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1436_ _1308_/X _1451_/A _1957_/B VGND VGND VPWR VPWR _1436_/Y sky130_fd_sc_hd__nor3_4
X_1505_ _1503_/X _1042_/A _1504_/X VGND VGND VPWR VPWR _1505_/X sky130_fd_sc_hd__o21a_4
X_1298_ _1052_/A _1085_/Y _1298_/C VGND VGND VPWR VPWR _1298_/Y sky130_fd_sc_hd__nand3_4
XFILLER_11_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1221_ _1221_/A VGND VGND VPWR VPWR _1708_/A sky130_fd_sc_hd__buf_2
XFILLER_6_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1152_ _1215_/A _1344_/C _1344_/D _1152_/D VGND VGND VPWR VPWR _1197_/A sky130_fd_sc_hd__nand4_4
X_1083_ _1147_/B VGND VGND VPWR VPWR _1125_/D sky130_fd_sc_hd__buf_2
XFILLER_45_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1985_ _1499_/B MISO_fromClient _1984_/Y VGND VGND VPWR VPWR MISO_toHost sky130_fd_sc_hd__o21a_4
XFILLER_20_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1419_ _1396_/A _1846_/A _1396_/C VGND VGND VPWR VPWR _1420_/C sky130_fd_sc_hd__nand3_4
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1770_ _1770_/A _1475_/A VGND VGND VPWR VPWR _1770_/Y sky130_fd_sc_hd__nand2_4
XFILLER_42_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1204_ _1182_/C _1152_/D VGND VGND VPWR VPWR _1344_/B sky130_fd_sc_hd__nor2_4
X_2184_ _2189_/CLK _2184_/D VGND VGND VPWR VPWR _1589_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1066_ _1064_/Y _1055_/A _1432_/C _1066_/D VGND VGND VPWR VPWR _1282_/B sky130_fd_sc_hd__nand4_4
X_1135_ _1070_/X _1126_/B _1098_/X VGND VGND VPWR VPWR _1135_/X sky130_fd_sc_hd__a21o_4
X_1968_ _1036_/B _2014_/Q _1694_/X _1449_/Y VGND VGND VPWR VPWR _1968_/X sky130_fd_sc_hd__a211o_4
X_1899_ _1899_/A _1899_/B _2001_/D VGND VGND VPWR VPWR _1899_/Y sky130_fd_sc_hd__nand3_4
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1822_ _2120_/Q _1822_/B VGND VGND VPWR VPWR _1822_/X sky130_fd_sc_hd__xor2_4
X_1753_ _1958_/A _1445_/A _1112_/A VGND VGND VPWR VPWR _1753_/Y sky130_fd_sc_hd__nand3_4
X_1684_ _1681_/A VGND VGND VPWR VPWR _1697_/A sky130_fd_sc_hd__buf_2
X_2167_ _2189_/CLK _1673_/X VGND VGND VPWR VPWR _2167_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2236_ _2228_/CLK _1122_/Y VGND VGND VPWR VPWR _2236_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1049_ _1049_/A VGND VGND VPWR VPWR _1049_/X sky130_fd_sc_hd__buf_2
X_1118_ _1109_/A _1116_/X _1117_/Y VGND VGND VPWR VPWR _1118_/Y sky130_fd_sc_hd__o21ai_4
X_2098_ _2091_/CLK _2098_/D VGND VGND VPWR VPWR _2098_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2021_ _2108_/CLK _1997_/Q VGND VGND VPWR VPWR DATA_TO_HASH[0] sky130_fd_sc_hd__dfxtp_4
XFILLER_50_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1805_ _2129_/Q _1804_/Y VGND VGND VPWR VPWR _1806_/A sky130_fd_sc_hd__xor2_4
X_1736_ _1734_/Y _1213_/A _1735_/Y VGND VGND VPWR VPWR _1736_/Y sky130_fd_sc_hd__a21oi_4
X_1598_ _1598_/A VGND VGND VPWR VPWR _1598_/Y sky130_fd_sc_hd__inv_2
X_1667_ _1660_/Y _1641_/X _1666_/Y VGND VGND VPWR VPWR _1667_/Y sky130_fd_sc_hd__a21oi_4
X_2219_ _2231_/CLK _2219_/D VGND VGND VPWR VPWR _2219_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1452_ _1450_/X _1480_/A _1293_/X VGND VGND VPWR VPWR _1452_/Y sky130_fd_sc_hd__a21oi_4
X_1521_ _1625_/A VGND VGND VPWR VPWR _1521_/X sky130_fd_sc_hd__buf_2
X_1383_ _1383_/A VGND VGND VPWR VPWR _1383_/Y sky130_fd_sc_hd__inv_2
X_2004_ _2189_/CLK _2004_/D VGND VGND VPWR VPWR _2028_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_50_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_7_0_addressalyzerBlock.SPI_CLK clkbuf_4_7_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2058_/CLK sky130_fd_sc_hd__clkbuf_1
X_1719_ _1483_/B VGND VGND VPWR VPWR _1719_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1504_ _1625_/A VGND VGND VPWR VPWR _1504_/X sky130_fd_sc_hd__buf_2
X_1366_ _1366_/A VGND VGND VPWR VPWR _1396_/A sky130_fd_sc_hd__inv_2
X_1435_ _1448_/A VGND VGND VPWR VPWR _1957_/B sky130_fd_sc_hd__inv_2
X_1297_ _1296_/Y _1282_/A _1282_/B _1282_/C _1085_/Y VGND VGND VPWR VPWR _1297_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_36_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1220_ _1344_/B _1344_/C _1344_/D VGND VGND VPWR VPWR _1221_/A sky130_fd_sc_hd__and3_4
X_1151_ _1184_/A VGND VGND VPWR VPWR _1152_/D sky130_fd_sc_hd__inv_2
XFILLER_45_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1082_ _1077_/Y _1080_/Y _1081_/Y VGND VGND VPWR VPWR _1082_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_60_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1984_ _1984_/A _1499_/B VGND VGND VPWR VPWR _1984_/Y sky130_fd_sc_hd__nand2_4
X_1418_ _1403_/Y _1416_/Y _1417_/X VGND VGND VPWR VPWR _1420_/A sky130_fd_sc_hd__o21ai_4
X_1349_ _1355_/A _1348_/Y VGND VGND VPWR VPWR _1349_/Y sky130_fd_sc_hd__nor2_4
XFILLER_51_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1203_ _1202_/Y _1362_/A VGND VGND VPWR VPWR _1203_/Y sky130_fd_sc_hd__nor2_4
X_2183_ _2189_/CLK _2183_/D VGND VGND VPWR VPWR _1589_/A sky130_fd_sc_hd__dfxtp_4
X_1134_ _1133_/X _1123_/X _1079_/X VGND VGND VPWR VPWR _1134_/Y sky130_fd_sc_hd__a21oi_4
X_1065_ _1065_/A VGND VGND VPWR VPWR _1432_/C sky130_fd_sc_hd__inv_2
X_1967_ _1282_/C _1966_/Y _1446_/X VGND VGND VPWR VPWR _2011_/D sky130_fd_sc_hd__a21oi_4
X_1898_ _1898_/A VGND VGND VPWR VPWR _1899_/A sky130_fd_sc_hd__inv_2
XFILLER_56_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1821_ _1825_/A _1821_/B _1826_/A _1825_/B VGND VGND VPWR VPWR _1822_/B sky130_fd_sc_hd__and4_4
X_1752_ _1739_/X _1748_/Y _1751_/Y VGND VGND VPWR VPWR _1752_/Y sky130_fd_sc_hd__o21ai_4
X_1683_ _1701_/A _2160_/Q VGND VGND VPWR VPWR _1683_/X sky130_fd_sc_hd__and2_4
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2166_ _2124_/CLK _2166_/D VGND VGND VPWR VPWR _2166_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1117_ _1109_/A _1106_/X _1116_/B _1108_/X _1957_/C VGND VGND VPWR VPWR _1117_/Y
+ sky130_fd_sc_hd__a41oi_4
X_2235_ _2228_/CLK _2235_/D VGND VGND VPWR VPWR _2235_/Q sky130_fd_sc_hd__dfxtp_4
X_2097_ _2137_/CLK _1875_/Y VGND VGND VPWR VPWR _2041_/D sky130_fd_sc_hd__dfxtp_4
X_1048_ _1182_/C _1310_/A _1311_/A _1048_/D VGND VGND VPWR VPWR _1049_/A sky130_fd_sc_hd__nand4_4
XFILLER_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2020_ _2171_/CLK _1767_/C VGND VGND VPWR VPWR _2019_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_62_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1804_ _2128_/Q _1810_/B _1376_/A _1810_/A VGND VGND VPWR VPWR _1804_/Y sky130_fd_sc_hd__nand4_4
X_1735_ _1213_/A _2141_/Q VGND VGND VPWR VPWR _1735_/Y sky130_fd_sc_hd__nor2_4
X_1666_ _1660_/Y _1641_/X _1969_/A VGND VGND VPWR VPWR _1666_/Y sky130_fd_sc_hd__o21ai_4
X_1597_ _1591_/Y _1675_/B _1596_/Y VGND VGND VPWR VPWR _1598_/A sky130_fd_sc_hd__nand3_4
XFILLER_53_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2149_ _2194_/CLK _1700_/X VGND VGND VPWR VPWR _2149_/Q sky130_fd_sc_hd__dfxtp_4
X_2218_ _2218_/CLK _1434_/Y VGND VGND VPWR VPWR _1426_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_30_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_m1_clk_local clkbuf_0_m1_clk_local/X VGND VGND VPWR VPWR clkbuf_2_3_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
X_1520_ _1501_/Y _2197_/Q _1519_/X VGND VGND VPWR VPWR _2205_/D sky130_fd_sc_hd__o21a_4
Xclkbuf_4_12_0_addressalyzerBlock.SPI_CLK clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2216_/CLK sky130_fd_sc_hd__clkbuf_1
X_1451_ _1451_/A _1451_/B _1451_/C VGND VGND VPWR VPWR _1451_/Y sky130_fd_sc_hd__nor3_4
X_1382_ _1857_/A _1154_/X _1166_/X _1381_/Y VGND VGND VPWR VPWR _1382_/X sky130_fd_sc_hd__a211o_4
XFILLER_35_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2003_ _2029_/CLK _1236_/A VGND VGND VPWR VPWR _2027_/D sky130_fd_sc_hd__dfxtp_4
X_1649_ _1649_/A _1648_/X _1649_/C _1649_/D VGND VGND VPWR VPWR _1649_/X sky130_fd_sc_hd__and4_4
X_1718_ _1714_/Y _1718_/B VGND VGND VPWR VPWR _1718_/Y sky130_fd_sc_hd__nand2_4
XFILLER_58_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1503_ _2215_/Q VGND VGND VPWR VPWR _1503_/X sky130_fd_sc_hd__buf_2
X_1365_ _1270_/Y VGND VGND VPWR VPWR _1397_/B sky130_fd_sc_hd__buf_2
X_1296_ _1086_/X _1049_/X _1110_/A VGND VGND VPWR VPWR _1296_/Y sky130_fd_sc_hd__o21ai_4
X_1434_ _1426_/Y _1430_/Y _1433_/X VGND VGND VPWR VPWR _1434_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_23_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1150_ _1182_/B VGND VGND VPWR VPWR _1344_/D sky130_fd_sc_hd__buf_2
Xclkbuf_3_4_0_m1_clk_local clkbuf_3_4_0_m1_clk_local/A VGND VGND VPWR VPWR _2108_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1081_ _1059_/B _1069_/B _1031_/X VGND VGND VPWR VPWR _1081_/Y sky130_fd_sc_hd__o21ai_4
X_1983_ _1983_/A VGND VGND VPWR VPWR _1984_/A sky130_fd_sc_hd__inv_2
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1417_ _1312_/X _1826_/A _1313_/B _1366_/A VGND VGND VPWR VPWR _1417_/X sky130_fd_sc_hd__a211o_4
X_1279_ _1278_/Y VGND VGND VPWR VPWR _1279_/Y sky130_fd_sc_hd__inv_2
X_1348_ _1348_/A VGND VGND VPWR VPWR _1348_/Y sky130_fd_sc_hd__inv_2
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1202_ _1202_/A VGND VGND VPWR VPWR _1202_/Y sky130_fd_sc_hd__inv_2
X_2182_ _2182_/CLK _1614_/Y VGND VGND VPWR VPWR _1574_/A sky130_fd_sc_hd__dfxtp_4
X_1064_ _1064_/A VGND VGND VPWR VPWR _1064_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1133_ _1904_/A VGND VGND VPWR VPWR _1133_/X sky130_fd_sc_hd__buf_2
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1966_ _1036_/B _1078_/X VGND VGND VPWR VPWR _1966_/Y sky130_fd_sc_hd__nand2_4
XFILLER_18_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1897_ _1217_/X _1896_/Y _1329_/X VGND VGND VPWR VPWR _1898_/A sky130_fd_sc_hd__and3_4
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1820_ _1820_/A _1819_/Y VGND VGND VPWR VPWR _1820_/X sky130_fd_sc_hd__xor2_4
XFILLER_47_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1751_ _1754_/A _1754_/B _1253_/A VGND VGND VPWR VPWR _1751_/Y sky130_fd_sc_hd__nand3_4
X_1682_ _1701_/A _2152_/Q VGND VGND VPWR VPWR _1682_/X sky130_fd_sc_hd__and2_4
XFILLER_38_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2234_ _2228_/CLK _1136_/Y VGND VGND VPWR VPWR _1108_/A sky130_fd_sc_hd__dfxtp_4
X_2165_ _2189_/CLK _1677_/X VGND VGND VPWR VPWR _1581_/B sky130_fd_sc_hd__dfxtp_4
X_1047_ _1047_/A VGND VGND VPWR VPWR _1311_/A sky130_fd_sc_hd__buf_2
X_1116_ _1052_/X _1116_/B _1108_/X _1125_/A VGND VGND VPWR VPWR _1116_/X sky130_fd_sc_hd__and4_4
X_2096_ _2137_/CLK _2096_/D VGND VGND VPWR VPWR _2040_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_21_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1949_ _1948_/X VGND VGND VPWR VPWR _1949_/X sky130_fd_sc_hd__buf_2
XFILLER_56_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1803_ _1803_/A _1787_/Y VGND VGND VPWR VPWR _1810_/B sky130_fd_sc_hd__nor2_4
X_1596_ _1600_/C _1596_/B _2185_/Q CLK_LED VGND VGND VPWR VPWR _1596_/Y sky130_fd_sc_hd__nand4_4
X_1734_ _1709_/X _1731_/Y _1733_/X VGND VGND VPWR VPWR _1734_/Y sky130_fd_sc_hd__o21ai_4
X_1665_ _1917_/A VGND VGND VPWR VPWR _1969_/A sky130_fd_sc_hd__buf_2
XFILLER_58_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2217_ _2248_/CLK _2217_/D VGND VGND VPWR VPWR _2217_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2079_ _2231_/CLK _1923_/Y VGND VGND VPWR VPWR _1773_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_41_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2148_ _2248_/CLK _1701_/Y VGND VGND VPWR VPWR _2148_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_30_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1450_ _1448_/A _1092_/A _1448_/Y _1449_/Y VGND VGND VPWR VPWR _1450_/X sky130_fd_sc_hd__a211o_4
X_1381_ _1355_/A _1380_/Y VGND VGND VPWR VPWR _1381_/Y sky130_fd_sc_hd__nor2_4
XFILLER_35_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2002_ _2182_/CLK _1258_/A VGND VGND VPWR VPWR _2026_/D sky130_fd_sc_hd__dfxtp_4
X_1648_ _1648_/A VGND VGND VPWR VPWR _1648_/X sky130_fd_sc_hd__buf_2
X_1579_ _1643_/A VGND VGND VPWR VPWR _1579_/Y sky130_fd_sc_hd__inv_2
X_1717_ _1715_/Y _1170_/X _1716_/Y VGND VGND VPWR VPWR _1718_/B sky130_fd_sc_hd__o21ai_4
XFILLER_58_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1433_ _1429_/X _1432_/Y _1293_/X VGND VGND VPWR VPWR _1433_/X sky130_fd_sc_hd__a21o_4
X_1502_ _1501_/Y VGND VGND VPWR VPWR _1573_/B sky130_fd_sc_hd__buf_2
X_1364_ _1346_/X _1361_/Y _1363_/X VGND VGND VPWR VPWR _1364_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_48_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1295_ _1289_/Y _1290_/Y _1294_/X VGND VGND VPWR VPWR _2228_/D sky130_fd_sc_hd__a21oi_4
XFILLER_23_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_addressalyzerBlock.SPI_CLK clkbuf_2_3_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1080_ _1892_/A _1078_/X _1079_/X VGND VGND VPWR VPWR _1080_/Y sky130_fd_sc_hd__a21oi_4
X_1982_ _1980_/Y S1_CLK_SELECT _1981_/Y VGND VGND VPWR VPWR _1982_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1416_ _1414_/Y _1285_/X _1415_/Y VGND VGND VPWR VPWR _1416_/Y sky130_fd_sc_hd__a21oi_4
X_1347_ _2142_/Q VGND VGND VPWR VPWR _1355_/A sky130_fd_sc_hd__buf_2
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1278_ _1064_/A _2012_/Q VGND VGND VPWR VPWR _1278_/Y sky130_fd_sc_hd__nor2_4
XFILLER_28_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1201_ _1311_/A _1201_/B VGND VGND VPWR VPWR _1202_/A sky130_fd_sc_hd__nor2_4
XFILLER_2_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1132_ _1108_/X _1106_/X _1129_/Y VGND VGND VPWR VPWR _1132_/Y sky130_fd_sc_hd__o21ai_4
X_2181_ _2182_/CLK _2181_/D VGND VGND VPWR VPWR _2181_/Q sky130_fd_sc_hd__dfxtp_4
X_1063_ _1092_/A _1066_/D _1280_/A VGND VGND VPWR VPWR _1282_/A sky130_fd_sc_hd__a21o_4
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1965_ _1964_/Y _1444_/Y _1446_/X VGND VGND VPWR VPWR _1965_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1896_ _1038_/A _1886_/C VGND VGND VPWR VPWR _1896_/Y sky130_fd_sc_hd__nor2_4
XFILLER_56_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1750_ _1008_/A VGND VGND VPWR VPWR _1754_/B sky130_fd_sc_hd__buf_2
XFILLER_15_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1681_ _1681_/A VGND VGND VPWR VPWR _1701_/A sky130_fd_sc_hd__buf_2
X_2164_ _2124_/CLK _2164_/D VGND VGND VPWR VPWR _1668_/A sky130_fd_sc_hd__dfxtp_4
X_2233_ _2051_/CLK _1142_/Y VGND VGND VPWR VPWR _1105_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1115_ _1678_/A _1115_/B VGND VGND VPWR VPWR _2237_/D sky130_fd_sc_hd__nor2_4
X_1046_ _1184_/A VGND VGND VPWR VPWR _1310_/A sky130_fd_sc_hd__buf_2
X_2095_ _2137_/CLK _1880_/Y VGND VGND VPWR VPWR _2039_/D sky130_fd_sc_hd__dfxtp_4
X_1879_ _1871_/X _1899_/B _2039_/D VGND VGND VPWR VPWR _1879_/Y sky130_fd_sc_hd__nand3_4
X_1948_ _1219_/B _1144_/B _1310_/X _1442_/X _1330_/A VGND VGND VPWR VPWR _1948_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1802_ _1790_/A _1802_/B VGND VGND VPWR VPWR _2130_/D sky130_fd_sc_hd__xnor2_4
X_1733_ _1215_/A _2043_/Q _1215_/B _1733_/D VGND VGND VPWR VPWR _1733_/X sky130_fd_sc_hd__or4_4
X_1595_ _1595_/A _1595_/B _1604_/A VGND VGND VPWR VPWR _1596_/B sky130_fd_sc_hd__nor3_4
X_1664_ _1664_/A VGND VGND VPWR VPWR _2169_/D sky130_fd_sc_hd__inv_2
X_2216_ _2216_/CLK _1454_/Y VGND VGND VPWR VPWR _1213_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_38_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2147_ _2218_/CLK _1702_/Y VGND VGND VPWR VPWR _2147_/Q sky130_fd_sc_hd__dfxtp_4
X_1029_ _2242_/Q _0998_/B _1028_/X VGND VGND VPWR VPWR _1029_/Y sky130_fd_sc_hd__o21ai_4
X_2078_ _2218_/CLK _1925_/Y VGND VGND VPWR VPWR _2078_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1380_ _2071_/Q VGND VGND VPWR VPWR _1380_/Y sky130_fd_sc_hd__inv_2
X_2001_ _2025_/CLK _2001_/D VGND VGND VPWR VPWR _2001_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_50_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1716_ _1170_/A _2037_/D _2143_/Q VGND VGND VPWR VPWR _1716_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_58_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1578_ _1648_/A VGND VGND VPWR VPWR _1578_/Y sky130_fd_sc_hd__inv_2
X_1647_ _1642_/B _1641_/X VGND VGND VPWR VPWR _1649_/A sky130_fd_sc_hd__nor2_4
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1363_ _1312_/X _2120_/Q _1313_/B _1366_/A VGND VGND VPWR VPWR _1363_/X sky130_fd_sc_hd__a211o_4
X_1432_ _1971_/A _1971_/C _1432_/C VGND VGND VPWR VPWR _1432_/Y sky130_fd_sc_hd__nand3_4
X_1501_ _2215_/Q VGND VGND VPWR VPWR _1501_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1294_ _1291_/X _1084_/Y _1293_/X VGND VGND VPWR VPWR _1294_/X sky130_fd_sc_hd__a21o_4
XFILLER_11_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1981_ _2192_/Q S1_CLK_SELECT VGND VGND VPWR VPWR _1981_/Y sky130_fd_sc_hd__nor2_4
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1346_ _1186_/Y _2128_/Q _1153_/Y VGND VGND VPWR VPWR _1346_/X sky130_fd_sc_hd__a21o_4
X_1415_ _1179_/X _2046_/Q _1187_/Y VGND VGND VPWR VPWR _1415_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_28_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1277_ _1089_/X _1087_/Y _1276_/Y VGND VGND VPWR VPWR _1277_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_59_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1200_ _1153_/Y _1193_/Y _1199_/X VGND VGND VPWR VPWR _1200_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_33_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2180_ _2182_/CLK _1623_/X VGND VGND VPWR VPWR _1587_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_2_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1062_ _1042_/Y _1066_/D _1061_/Y VGND VGND VPWR VPWR _1062_/Y sky130_fd_sc_hd__o21ai_4
X_1131_ _1128_/Y _1130_/Y _1040_/X VGND VGND VPWR VPWR _2235_/D sky130_fd_sc_hd__a21oi_4
X_1964_ _1030_/X _2014_/Q VGND VGND VPWR VPWR _1964_/Y sky130_fd_sc_hd__nand2_4
X_1895_ _1894_/Y _1885_/X _1888_/X _1258_/Y _1890_/X VGND VGND VPWR VPWR _2090_/D
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_3_0_0_m1_clk_local clkbuf_3_1_0_m1_clk_local/A VGND VGND VPWR VPWR _2182_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_1329_ _1152_/D VGND VGND VPWR VPWR _1329_/X sky130_fd_sc_hd__buf_2
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1680_ _1678_/A _1693_/B VGND VGND VPWR VPWR _2163_/D sky130_fd_sc_hd__nor2_4
X_2232_ _2231_/CLK _2232_/D VGND VGND VPWR VPWR _1228_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_38_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1114_ _1057_/A _1111_/X _1113_/Y _1069_/B VGND VGND VPWR VPWR _1115_/B sky130_fd_sc_hd__a22oi_4
X_2163_ _2218_/CLK _2163_/D VGND VGND VPWR VPWR _1693_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1045_ _1149_/B VGND VGND VPWR VPWR _1086_/A sky130_fd_sc_hd__inv_2
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2094_ _2137_/CLK _2094_/D VGND VGND VPWR VPWR _2038_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_21_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1878_ _1756_/Y _1865_/X _1877_/Y VGND VGND VPWR VPWR _2096_/D sky130_fd_sc_hd__o21ai_4
XFILLER_9_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1947_ _1892_/Y _1943_/Y _1946_/Y VGND VGND VPWR VPWR _2067_/D sky130_fd_sc_hd__o21ai_4
XFILLER_56_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1801_ _2129_/Q _1797_/Y _1807_/A _1376_/A VGND VGND VPWR VPWR _1802_/B sky130_fd_sc_hd__nand4_4
X_1732_ _1243_/C VGND VGND VPWR VPWR _1733_/D sky130_fd_sc_hd__buf_2
X_1663_ _1580_/B _1661_/Y _1662_/Y VGND VGND VPWR VPWR _1664_/A sky130_fd_sc_hd__a21o_4
XFILLER_7_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1594_ _1588_/B VGND VGND VPWR VPWR _1604_/A sky130_fd_sc_hd__buf_2
XFILLER_38_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2077_ _2085_/CLK _1926_/Y VGND VGND VPWR VPWR _2017_/D sky130_fd_sc_hd__dfxtp_4
X_2215_ _2218_/CLK _2215_/D VGND VGND VPWR VPWR _2215_/Q sky130_fd_sc_hd__dfxtp_4
X_2146_ _2248_/CLK _2146_/D VGND VGND VPWR VPWR _2146_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1028_ _1034_/C _0996_/A VGND VGND VPWR VPWR _1028_/X sky130_fd_sc_hd__or2_4
XFILLER_34_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2000_ _2182_/CLK _2088_/Q VGND VGND VPWR VPWR _2024_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_50_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_3_0_addressalyzerBlock.SPI_CLK clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR clkbuf_4_7_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_23_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1646_ _1646_/A _1675_/B _1646_/C VGND VGND VPWR VPWR _2174_/D sky130_fd_sc_hd__and3_4
X_1715_ _1997_/D VGND VGND VPWR VPWR _1715_/Y sky130_fd_sc_hd__inv_2
X_1577_ _1609_/B VGND VGND VPWR VPWR _1584_/C sky130_fd_sc_hd__inv_2
X_2129_ _2124_/CLK _2129_/D VGND VGND VPWR VPWR _2129_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1500_ _1498_/Y _1499_/Y _1446_/X VGND VGND VPWR VPWR _1500_/Y sky130_fd_sc_hd__a21oi_4
X_1362_ _1362_/A VGND VGND VPWR VPWR _1366_/A sky130_fd_sc_hd__buf_2
X_1431_ _1431_/A VGND VGND VPWR VPWR _1971_/C sky130_fd_sc_hd__inv_2
X_1293_ _1330_/A VGND VGND VPWR VPWR _1293_/X sky130_fd_sc_hd__buf_2
XFILLER_51_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1629_ _1628_/Y VGND VGND VPWR VPWR _2179_/D sky130_fd_sc_hd__inv_2
XFILLER_54_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1980_ S1_CLK_IN VGND VGND VPWR VPWR _1980_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1345_ _1344_/X VGND VGND VPWR VPWR _1421_/A sky130_fd_sc_hd__buf_2
X_1276_ _1089_/X _1052_/A _1125_/D _1149_/A _1957_/C VGND VGND VPWR VPWR _1276_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1414_ _1410_/X _1413_/X VGND VGND VPWR VPWR _1414_/Y sky130_fd_sc_hd__nand2_4
XFILLER_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1130_ _1070_/X _1129_/Y _1116_/B VGND VGND VPWR VPWR _1130_/Y sky130_fd_sc_hd__o21ai_4
X_1061_ _1044_/Y _1053_/X _1110_/A _1061_/D VGND VGND VPWR VPWR _1061_/Y sky130_fd_sc_hd__nand4_4
XFILLER_18_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1963_ _1678_/A _1962_/Y VGND VGND VPWR VPWR _2012_/D sky130_fd_sc_hd__nor2_4
X_1894_ _1894_/A VGND VGND VPWR VPWR _1894_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1328_ _1310_/X _1207_/B _1314_/X VGND VGND VPWR VPWR _1328_/Y sky130_fd_sc_hd__o21ai_4
X_1259_ _1171_/X _2098_/Q _2143_/Q VGND VGND VPWR VPWR _1259_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2231_ _2231_/CLK _2231_/D VGND VGND VPWR VPWR _2231_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_2_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1044_ _2240_/Q VGND VGND VPWR VPWR _1044_/Y sky130_fd_sc_hd__inv_2
X_1113_ _1057_/A _1071_/X _1109_/Y _1112_/Y _1066_/D VGND VGND VPWR VPWR _1113_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_0_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2093_ _2211_/CLK _2093_/D VGND VGND VPWR VPWR _2037_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2162_ _2218_/CLK _1682_/X VGND VGND VPWR VPWR _1679_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_61_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1877_ _1871_/X _1899_/B _2040_/D VGND VGND VPWR VPWR _1877_/Y sky130_fd_sc_hd__nand3_4
X_1946_ _1943_/Y _1341_/C _1484_/B VGND VGND VPWR VPWR _1946_/Y sky130_fd_sc_hd__nand3_4
XFILLER_29_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1800_ _1800_/A VGND VGND VPWR VPWR _2131_/D sky130_fd_sc_hd__inv_2
XFILLER_34_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1731_ _1710_/Y _1730_/Y VGND VGND VPWR VPWR _1731_/Y sky130_fd_sc_hd__nor2_4
X_1662_ _1580_/B _1661_/Y _1681_/A VGND VGND VPWR VPWR _1662_/Y sky130_fd_sc_hd__o21ai_4
X_2214_ _2231_/CLK _1481_/X VGND VGND VPWR VPWR _1480_/B sky130_fd_sc_hd__dfxtp_4
X_1593_ _1589_/A VGND VGND VPWR VPWR _1595_/B sky130_fd_sc_hd__inv_2
X_1027_ _1025_/Y _1003_/X _1026_/Y VGND VGND VPWR VPWR _1027_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_26_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2145_ _2248_/CLK _2145_/D VGND VGND VPWR VPWR _1703_/B sky130_fd_sc_hd__dfxtp_4
X_2076_ _2091_/CLK _2076_/D VGND VGND VPWR VPWR _2076_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_19_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1929_ _1927_/Y _1341_/C _2076_/Q _1185_/A _1928_/Y VGND VGND VPWR VPWR _2076_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_39_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1645_ _1642_/Y _1649_/C _1649_/D _2173_/Q _2174_/Q VGND VGND VPWR VPWR _1646_/A
+ sky130_fd_sc_hd__a41o_4
X_1576_ _1576_/A VGND VGND VPWR VPWR _1584_/B sky130_fd_sc_hd__inv_2
X_1714_ _1712_/Y _1170_/X _1713_/Y VGND VGND VPWR VPWR _1714_/Y sky130_fd_sc_hd__o21ai_4
X_2128_ _2124_/CLK _1808_/Y VGND VGND VPWR VPWR _2128_/Q sky130_fd_sc_hd__dfxtp_4
X_2059_ _2044_/CLK DATA_FROM_HASH[6] VGND VGND VPWR VPWR _2059_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1430_ _1308_/X _1969_/D _1431_/A _1065_/A _1429_/X VGND VGND VPWR VPWR _1430_/Y
+ sky130_fd_sc_hd__o41ai_4
X_1361_ _1359_/Y _1285_/X _1360_/Y VGND VGND VPWR VPWR _1361_/Y sky130_fd_sc_hd__a21oi_4
X_1292_ _1038_/A VGND VGND VPWR VPWR _1330_/A sky130_fd_sc_hd__buf_2
XFILLER_63_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1559_ _2192_/Q _1565_/A SPI_CLK_RESET_N VGND VGND VPWR VPWR _1559_/Y sky130_fd_sc_hd__o21ai_4
X_1628_ _1628_/A _1628_/B VGND VGND VPWR VPWR _1628_/Y sky130_fd_sc_hd__nand2_4
XFILLER_36_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1413_ _1763_/C _1355_/X _1161_/A _1412_/Y VGND VGND VPWR VPWR _1413_/X sky130_fd_sc_hd__a211o_4
X_1275_ _1275_/A _1275_/B VGND VGND VPWR VPWR _1275_/Y sky130_fd_sc_hd__nand2_4
X_1344_ _1344_/A _1344_/B _1344_/C _1344_/D VGND VGND VPWR VPWR _1344_/X sky130_fd_sc_hd__and4_4
XFILLER_3_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1060_ _1059_/X VGND VGND VPWR VPWR _1061_/D sky130_fd_sc_hd__buf_2
XFILLER_33_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1962_ _2158_/Q _1065_/A _1030_/X _1078_/X VGND VGND VPWR VPWR _1962_/Y sky130_fd_sc_hd__a22oi_4
X_1893_ _1892_/Y _1885_/X _1888_/X _1236_/Y _1890_/X VGND VGND VPWR VPWR _2091_/D
+ sky130_fd_sc_hd__o32ai_4
X_1189_ _1189_/A VGND VGND VPWR VPWR _1243_/B sky130_fd_sc_hd__buf_2
XFILLER_24_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1258_ _1258_/A VGND VGND VPWR VPWR _1258_/Y sky130_fd_sc_hd__inv_2
X_1327_ _1969_/D _1123_/X _1902_/A VGND VGND VPWR VPWR _1327_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_33_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2230_ _2052_/CLK _1275_/Y VGND VGND VPWR VPWR _2230_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2161_ _2248_/CLK _1683_/X VGND VGND VPWR VPWR _2161_/Q sky130_fd_sc_hd__dfxtp_4
X_1043_ _2012_/Q VGND VGND VPWR VPWR _1066_/D sky130_fd_sc_hd__inv_2
X_1112_ _1112_/A VGND VGND VPWR VPWR _1112_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2092_ _2085_/CLK _1891_/Y VGND VGND VPWR VPWR _2004_/D sky130_fd_sc_hd__dfxtp_4
X_1945_ _1042_/Y _1943_/Y _1944_/Y VGND VGND VPWR VPWR _2068_/D sky130_fd_sc_hd__o21ai_4
X_1876_ _1008_/A VGND VGND VPWR VPWR _1899_/B sky130_fd_sc_hd__buf_2
XFILLER_56_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_3_0_addressalyzerBlock.SPI_CLK clkbuf_4_3_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2224_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_62_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1730_ _1725_/Y _1727_/X _1729_/Y VGND VGND VPWR VPWR _1730_/Y sky130_fd_sc_hd__a21oi_4
X_1592_ _1589_/C VGND VGND VPWR VPWR _1600_/C sky130_fd_sc_hd__buf_2
X_1661_ _1660_/Y _1641_/X VGND VGND VPWR VPWR _1661_/Y sky130_fd_sc_hd__nor2_4
XFILLER_11_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2144_ _2224_/CLK _2144_/D VGND VGND VPWR VPWR _2144_/Q sky130_fd_sc_hd__dfxtp_4
X_2213_ _2213_/CLK _2213_/D VGND VGND VPWR VPWR _2213_/Q sky130_fd_sc_hd__dfxtp_4
X_1026_ _1400_/B _1003_/A _1008_/X VGND VGND VPWR VPWR _1026_/Y sky130_fd_sc_hd__o21ai_4
X_2075_ _2091_/CLK _2075_/D VGND VGND VPWR VPWR _2075_/Q sky130_fd_sc_hd__dfxtp_4
X_1859_ _1858_/X VGND VGND VPWR VPWR _2103_/D sky130_fd_sc_hd__inv_2
X_1928_ _1741_/Y VGND VGND VPWR VPWR _1928_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_2_2_0_m1_clk_local clkbuf_2_3_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_3_4_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1713_ _1171_/X _2030_/D _1166_/A VGND VGND VPWR VPWR _1713_/Y sky130_fd_sc_hd__a21oi_4
X_1644_ _1583_/A VGND VGND VPWR VPWR _1649_/D sky130_fd_sc_hd__buf_2
X_1575_ _2175_/Q VGND VGND VPWR VPWR _1575_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2127_ _2124_/CLK _2127_/D VGND VGND VPWR VPWR _1376_/A sky130_fd_sc_hd__dfxtp_4
X_2058_ _2058_/CLK DATA_FROM_HASH[5] VGND VGND VPWR VPWR _2050_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_41_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1009_ _2231_/Q _1004_/X _1008_/X VGND VGND VPWR VPWR _1009_/Y sky130_fd_sc_hd__o21ai_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1360_ _1285_/X _2048_/Q _1188_/X VGND VGND VPWR VPWR _1360_/Y sky130_fd_sc_hd__o21ai_4
X_1291_ _1291_/A VGND VGND VPWR VPWR _1291_/X sky130_fd_sc_hd__buf_2
XFILLER_36_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1558_ _1563_/A _1562_/C _1570_/C VGND VGND VPWR VPWR _1565_/A sky130_fd_sc_hd__nor3_4
X_1489_ _1487_/Y _1057_/A _1109_/A _1356_/Y VGND VGND VPWR VPWR _1489_/Y sky130_fd_sc_hd__a22oi_4
X_1627_ _1621_/C _1608_/Y _1624_/D _1627_/D VGND VGND VPWR VPWR _1628_/B sky130_fd_sc_hd__nand4_4
XFILLER_10_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1343_ _1217_/X _1708_/A _1480_/A _1215_/Y VGND VGND VPWR VPWR _1343_/X sky130_fd_sc_hd__a211o_4
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1412_ _1412_/A _1411_/Y VGND VGND VPWR VPWR _1412_/Y sky130_fd_sc_hd__nor2_4
X_1274_ _1274_/A _2230_/Q VGND VGND VPWR VPWR _1275_/B sky130_fd_sc_hd__nand2_4
XFILLER_36_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1961_ _1656_/A _1030_/X _1971_/C _1971_/B _1960_/X VGND VGND VPWR VPWR _2008_/D
+ sky130_fd_sc_hd__o32ai_4
X_1892_ _1892_/A VGND VGND VPWR VPWR _1892_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1326_ _1326_/A VGND VGND VPWR VPWR _1902_/A sky130_fd_sc_hd__buf_2
X_1188_ _1187_/Y VGND VGND VPWR VPWR _1188_/X sky130_fd_sc_hd__buf_2
XFILLER_24_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1257_ _1255_/Y _1233_/X _1256_/Y VGND VGND VPWR VPWR _1257_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_59_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE2_0 _1236_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2160_ _2194_/CLK _1685_/X VGND VGND VPWR VPWR _2160_/Q sky130_fd_sc_hd__dfxtp_4
X_1111_ _1109_/Y _1298_/C _1067_/Y VGND VGND VPWR VPWR _1111_/X sky130_fd_sc_hd__a21o_4
X_1042_ _1042_/A VGND VGND VPWR VPWR _1042_/Y sky130_fd_sc_hd__inv_2
X_2091_ _2091_/CLK _2091_/D VGND VGND VPWR VPWR _1236_/A sky130_fd_sc_hd__dfxtp_4
X_1875_ _1753_/Y _1865_/X _1874_/Y VGND VGND VPWR VPWR _1875_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_14_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1944_ _1943_/Y _1917_/X _1944_/C VGND VGND VPWR VPWR _1944_/Y sky130_fd_sc_hd__nand3_4
XFILLER_21_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1309_ _1449_/B VGND VGND VPWR VPWR _1451_/A sky130_fd_sc_hd__buf_2
XFILLER_28_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1591_ _1589_/Y _1591_/B VGND VGND VPWR VPWR _1591_/Y sky130_fd_sc_hd__nand2_4
X_1660_ _2168_/Q VGND VGND VPWR VPWR _1660_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2143_ _2051_/CLK _2143_/D VGND VGND VPWR VPWR _2143_/Q sky130_fd_sc_hd__dfxtp_4
X_2212_ _2218_/CLK _1500_/Y VGND VGND VPWR VPWR _1499_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1025_ _2242_/Q _0996_/A _1024_/X VGND VGND VPWR VPWR _1025_/Y sky130_fd_sc_hd__o21ai_4
X_2074_ _2091_/CLK _2074_/D VGND VGND VPWR VPWR _2074_/Q sky130_fd_sc_hd__dfxtp_4
X_1858_ _1773_/B _1858_/B VGND VGND VPWR VPWR _1858_/X sky130_fd_sc_hd__xor2_4
X_1927_ _1329_/X _1144_/B _1196_/X _1442_/X VGND VGND VPWR VPWR _1927_/Y sky130_fd_sc_hd__nand4_4
X_1789_ _2128_/Q VGND VGND VPWR VPWR _1807_/A sky130_fd_sc_hd__buf_2
XFILLER_39_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1643_ _1643_/A VGND VGND VPWR VPWR _1649_/C sky130_fd_sc_hd__buf_2
XFILLER_31_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1712_ _2017_/D VGND VGND VPWR VPWR _1712_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1574_ _1574_/A VGND VGND VPWR VPWR _1595_/A sky130_fd_sc_hd__inv_2
XFILLER_6_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2126_ _2124_/CLK _2126_/D VGND VGND VPWR VPWR _1810_/A sky130_fd_sc_hd__dfxtp_4
X_2057_ _2211_/CLK DATA_FROM_HASH[4] VGND VGND VPWR VPWR _2049_/D sky130_fd_sc_hd__dfxtp_4
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1008_ _1008_/A VGND VGND VPWR VPWR _1008_/X sky130_fd_sc_hd__buf_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1290_ _1892_/A _1279_/Y _1306_/A VGND VGND VPWR VPWR _1290_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_31_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1626_ _1627_/D _1624_/X _1681_/A VGND VGND VPWR VPWR _1628_/A sky130_fd_sc_hd__o21a_4
X_1557_ _1569_/A _2189_/Q VGND VGND VPWR VPWR _1570_/C sky130_fd_sc_hd__nand2_4
XFILLER_39_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1488_ _1057_/A _1487_/Y _2235_/Q _1389_/B VGND VGND VPWR VPWR _1488_/X sky130_fd_sc_hd__o22a_4
X_2109_ _2115_/CLK _1848_/Y VGND VGND VPWR VPWR _2109_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1273_ _1268_/Y _1269_/Y _1272_/X VGND VGND VPWR VPWR _1275_/A sky130_fd_sc_hd__a21o_4
X_1342_ _1341_/Y VGND VGND VPWR VPWR _1342_/Y sky130_fd_sc_hd__inv_2
X_1411_ _1482_/A VGND VGND VPWR VPWR _1411_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1609_ _1608_/Y _1609_/B _1587_/A _1587_/D VGND VGND VPWR VPWR _1609_/X sky130_fd_sc_hd__and4_4
XFILLER_59_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1960_ _1003_/A _1972_/C _1330_/X VGND VGND VPWR VPWR _1960_/X sky130_fd_sc_hd__a21o_4
X_1891_ _1042_/Y _1885_/X _1888_/X _1169_/Y _1890_/X VGND VGND VPWR VPWR _1891_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1325_ _1064_/A VGND VGND VPWR VPWR _1969_/D sky130_fd_sc_hd__buf_2
X_1256_ _1164_/X _2074_/Q _1166_/A VGND VGND VPWR VPWR _1256_/Y sky130_fd_sc_hd__a21oi_4
X_1187_ _1186_/Y VGND VGND VPWR VPWR _1187_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_8_0_addressalyzerBlock.SPI_CLK clkbuf_4_9_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2211_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1110_ _1110_/A VGND VGND VPWR VPWR _1298_/C sky130_fd_sc_hd__buf_2
X_2090_ _2085_/CLK _2090_/D VGND VGND VPWR VPWR _1258_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1041_ _1034_/Y _1036_/Y _1040_/X VGND VGND VPWR VPWR _1041_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_21_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1874_ _1871_/X _1767_/B _2041_/D VGND VGND VPWR VPWR _1874_/Y sky130_fd_sc_hd__nand3_4
X_1943_ _1943_/A VGND VGND VPWR VPWR _1943_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1308_ _2010_/Q VGND VGND VPWR VPWR _1308_/X sky130_fd_sc_hd__buf_2
X_1239_ _1235_/Y _1238_/Y _1175_/X VGND VGND VPWR VPWR _1239_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1590_ CLK_LED VGND VGND VPWR VPWR _1591_/B sky130_fd_sc_hd__inv_2
XFILLER_53_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1024_ _1024_/A _1020_/B VGND VGND VPWR VPWR _1024_/X sky130_fd_sc_hd__or2_4
XFILLER_38_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2211_ _2211_/CLK _2211_/D VGND VGND VPWR VPWR _1042_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2073_ _2213_/CLK _1936_/Y VGND VGND VPWR VPWR _1462_/A sky130_fd_sc_hd__dfxtp_4
X_2142_ _2224_/CLK _2142_/D VGND VGND VPWR VPWR _2142_/Q sky130_fd_sc_hd__dfxtp_4
X_1788_ _1788_/A _1402_/Y _1803_/A _1787_/Y VGND VGND VPWR VPWR _1807_/B sky130_fd_sc_hd__nor4_4
X_1857_ _1857_/A _2102_/Q _2101_/Q VGND VGND VPWR VPWR _1858_/B sky130_fd_sc_hd__nand3_4
X_1926_ _1907_/Y _1909_/X _1887_/Y _1712_/Y _1910_/X VGND VGND VPWR VPWR _1926_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_55_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1711_ _1179_/X _2045_/Q _1187_/Y VGND VGND VPWR VPWR _1711_/Y sky130_fd_sc_hd__o21ai_4
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1642_ _1578_/Y _1642_/B _1641_/X VGND VGND VPWR VPWR _1642_/Y sky130_fd_sc_hd__nor3_4
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1573_ _1678_/A _1573_/B VGND VGND VPWR VPWR _1573_/Y sky130_fd_sc_hd__nor2_4
X_2125_ _2124_/CLK _2125_/D VGND VGND VPWR VPWR _1769_/A sky130_fd_sc_hd__dfxtp_4
X_2056_ _2211_/CLK DATA_FROM_HASH[3] VGND VGND VPWR VPWR _2056_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1007_ _1625_/A VGND VGND VPWR VPWR _1008_/A sky130_fd_sc_hd__buf_2
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1909_ _1206_/A VGND VGND VPWR VPWR _1909_/X sky130_fd_sc_hd__buf_2
XFILLER_57_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1556_ _0998_/B _1455_/D _1555_/Y VGND VGND VPWR VPWR _2193_/D sky130_fd_sc_hd__o21a_4
X_1625_ _1625_/A VGND VGND VPWR VPWR _1681_/A sky130_fd_sc_hd__buf_2
XFILLER_39_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1487_ _2065_/Q VGND VGND VPWR VPWR _1487_/Y sky130_fd_sc_hd__inv_2
X_2108_ _2108_/CLK _1850_/Y VGND VGND VPWR VPWR _1779_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_54_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2039_ _2182_/CLK _2039_/D VGND VGND VPWR VPWR _2033_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_10_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1410_ _1406_/X _1409_/Y _2144_/Q VGND VGND VPWR VPWR _1410_/X sky130_fd_sc_hd__a21o_4
X_1272_ _1271_/Y _1272_/B VGND VGND VPWR VPWR _1272_/X sky130_fd_sc_hd__or2_4
X_1341_ _1341_/A _1341_/B _1341_/C VGND VGND VPWR VPWR _1341_/Y sky130_fd_sc_hd__nand3_4
XFILLER_36_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1608_ _1607_/X _1584_/B _1583_/Y VGND VGND VPWR VPWR _1608_/Y sky130_fd_sc_hd__nor3_4
X_1539_ _2197_/Q _1524_/Y _1538_/X VGND VGND VPWR VPWR _2198_/D sky130_fd_sc_hd__o21a_4
XFILLER_47_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1890_ _1889_/X VGND VGND VPWR VPWR _1890_/X sky130_fd_sc_hd__buf_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1186_ _1189_/A _1185_/Y VGND VGND VPWR VPWR _1186_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_4_13_0_addressalyzerBlock.SPI_CLK clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2231_/CLK sky130_fd_sc_hd__clkbuf_1
X_1324_ _1315_/Y _1323_/Y _1040_/X VGND VGND VPWR VPWR _1324_/Y sky130_fd_sc_hd__a21oi_4
X_1255_ ID_toHost VGND VGND VPWR VPWR _1255_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_7_0_m1_clk_local clkbuf_3_7_0_m1_clk_local/A VGND VGND VPWR VPWR _2115_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1040_ _1040_/A VGND VGND VPWR VPWR _1040_/X sky130_fd_sc_hd__buf_2
XFILLER_64_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1942_ _1396_/C _1005_/Y _1310_/X _2217_/Q VGND VGND VPWR VPWR _1943_/A sky130_fd_sc_hd__and4_4
X_1873_ _1748_/Y _1865_/X _1872_/Y VGND VGND VPWR VPWR _2098_/D sky130_fd_sc_hd__o21ai_4
XFILLER_9_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1307_ _1307_/A _1675_/B _1307_/C VGND VGND VPWR VPWR _1307_/X sky130_fd_sc_hd__and3_4
X_1238_ _1236_/Y _1170_/X _1237_/Y VGND VGND VPWR VPWR _1238_/Y sky130_fd_sc_hd__o21ai_4
X_1169_ _2004_/D VGND VGND VPWR VPWR _1169_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2210_ _2211_/CLK _1508_/X VGND VGND VPWR VPWR _1892_/A sky130_fd_sc_hd__dfxtp_4
X_1023_ _1021_/Y _1003_/X _1022_/Y VGND VGND VPWR VPWR _2244_/D sky130_fd_sc_hd__a21oi_4
X_2141_ _2216_/CLK _1736_/Y VGND VGND VPWR VPWR _2141_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_34_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2072_ _2211_/CLK _2072_/D VGND VGND VPWR VPWR _1348_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_34_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1925_ _1904_/Y _1916_/X _1924_/Y VGND VGND VPWR VPWR _1925_/Y sky130_fd_sc_hd__o21ai_4
X_1787_ _1825_/A _1815_/B _1815_/C _1787_/D VGND VGND VPWR VPWR _1787_/Y sky130_fd_sc_hd__nand4_4
X_1856_ _1371_/X _1774_/D VGND VGND VPWR VPWR _1856_/X sky130_fd_sc_hd__xor2_4
XFILLER_52_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1572_ _1569_/A _1572_/B VGND VGND VPWR VPWR _2188_/D sky130_fd_sc_hd__nor2_4
X_1710_ _2101_/Q _1270_/Y _1421_/Y VGND VGND VPWR VPWR _1710_/Y sky130_fd_sc_hd__o21ai_4
X_1641_ _1581_/Y VGND VGND VPWR VPWR _1641_/X sky130_fd_sc_hd__buf_2
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2124_ _2124_/CLK _1814_/Y VGND VGND VPWR VPWR _2124_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_3_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2055_ _2058_/CLK DATA_FROM_HASH[2] VGND VGND VPWR VPWR _2047_/D sky130_fd_sc_hd__dfxtp_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1006_ _1005_/Y VGND VGND VPWR VPWR _1625_/A sky130_fd_sc_hd__buf_2
XFILLER_22_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1839_ _1770_/A _1839_/B VGND VGND VPWR VPWR _1839_/X sky130_fd_sc_hd__xor2_4
X_1908_ _1907_/Y _1473_/B _1905_/X _1715_/Y _1889_/X VGND VGND VPWR VPWR _1908_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_22_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1624_ _1619_/Y _1621_/B _1609_/B _1624_/D VGND VGND VPWR VPWR _1624_/X sky130_fd_sc_hd__and4_4
X_1555_ _1555_/A VGND VGND VPWR VPWR _1555_/Y sky130_fd_sc_hd__inv_2
X_2107_ _2115_/CLK _1851_/X VGND VGND VPWR VPWR _1834_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_54_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1486_ _1486_/A VGND VGND VPWR VPWR _1486_/Y sky130_fd_sc_hd__inv_2
X_2038_ _2124_/CLK _2038_/D VGND VGND VPWR VPWR _2038_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_60_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1340_ _1917_/A VGND VGND VPWR VPWR _1341_/C sky130_fd_sc_hd__buf_2
X_1271_ _1772_/A _1270_/Y VGND VGND VPWR VPWR _1271_/Y sky130_fd_sc_hd__nor2_4
XFILLER_36_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1469_ _1189_/A _1190_/X _1052_/B _2049_/Q VGND VGND VPWR VPWR _1469_/Y sky130_fd_sc_hd__a2bb2oi_4
X_1607_ _1575_/Y VGND VGND VPWR VPWR _1607_/X sky130_fd_sc_hd__buf_2
X_1538_ _2198_/Q _2156_/Q _1535_/X VGND VGND VPWR VPWR _1538_/X sky130_fd_sc_hd__o21a_4
XFILLER_42_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1323_ _1317_/Y _1318_/X _1323_/C VGND VGND VPWR VPWR _1323_/Y sky130_fd_sc_hd__nand3_4
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1185_ _1185_/A VGND VGND VPWR VPWR _1185_/Y sky130_fd_sc_hd__inv_2
X_1254_ _1159_/X _1490_/A _1161_/X VGND VGND VPWR VPWR _1254_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_32_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1941_ _1927_/Y _1958_/A _2030_/D _1185_/A _1940_/Y VGND VGND VPWR VPWR _1941_/X
+ sky130_fd_sc_hd__a32o_4
X_1872_ _1871_/X _1767_/B _2098_/Q VGND VGND VPWR VPWR _1872_/Y sky130_fd_sc_hd__nand3_4
XFILLER_14_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1306_ _1306_/A _1086_/X VGND VGND VPWR VPWR _1307_/C sky130_fd_sc_hd__nand2_4
XFILLER_64_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1099_ _1070_/X _1097_/Y _1098_/X VGND VGND VPWR VPWR _1099_/X sky130_fd_sc_hd__a21o_4
X_1237_ _1171_/X _1869_/C _2143_/Q VGND VGND VPWR VPWR _1237_/Y sky130_fd_sc_hd__a21oi_4
X_1168_ _1163_/Y _1159_/X _1167_/Y VGND VGND VPWR VPWR _1168_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2140_ _2137_/CLK _2140_/D VGND VGND VPWR VPWR _1156_/A sky130_fd_sc_hd__dfxtp_4
X_1022_ _1374_/B _1004_/X _1008_/X VGND VGND VPWR VPWR _1022_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_38_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2071_ _2213_/CLK _1938_/Y VGND VGND VPWR VPWR _2071_/Q sky130_fd_sc_hd__dfxtp_4
X_1855_ _2105_/Q _1854_/Y VGND VGND VPWR VPWR _1855_/X sky130_fd_sc_hd__xor2_4
X_1924_ _1915_/Y _1917_/X _2078_/Q VGND VGND VPWR VPWR _1924_/Y sky130_fd_sc_hd__nand3_4
X_1786_ _1785_/Y VGND VGND VPWR VPWR _1787_/D sky130_fd_sc_hd__inv_2
XFILLER_37_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1571_ SPI_CLK_RESET_N VGND VGND VPWR VPWR _1572_/B sky130_fd_sc_hd__inv_2
X_1640_ _1607_/X _1646_/C _1639_/Y VGND VGND VPWR VPWR _1640_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2123_ _2025_/CLK _2123_/D VGND VGND VPWR VPWR _1813_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_54_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2054_ _2044_/CLK DATA_FROM_HASH[1] VGND VGND VPWR VPWR _2046_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_34_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1005_ _2006_/Q VGND VGND VPWR VPWR _1005_/Y sky130_fd_sc_hd__inv_2
X_1838_ _1840_/A _1840_/B VGND VGND VPWR VPWR _1839_/B sky130_fd_sc_hd__nor2_4
X_1907_ _1907_/A VGND VGND VPWR VPWR _1907_/Y sky130_fd_sc_hd__inv_2
X_1769_ _1769_/A VGND VGND VPWR VPWR _1803_/A sky130_fd_sc_hd__inv_2
XFILLER_25_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1623_ _1587_/A _1621_/X _1622_/Y VGND VGND VPWR VPWR _1623_/X sky130_fd_sc_hd__o21a_4
X_1485_ _1097_/Y _1490_/A _1482_/Y _1483_/X _1484_/X VGND VGND VPWR VPWR _1486_/A
+ sky130_fd_sc_hd__a2111o_4
X_1554_ _1549_/A _1535_/X _1553_/Y VGND VGND VPWR VPWR _1555_/A sky130_fd_sc_hd__nand3_4
.ends

