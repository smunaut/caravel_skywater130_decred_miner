VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 87.460 2924.800 88.660 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1984.510 2429.200 1984.830 2429.260 ;
        RECT 2898.070 2429.200 2898.390 2429.260 ;
        RECT 1984.510 2429.060 2898.390 2429.200 ;
        RECT 1984.510 2429.000 1984.830 2429.060 ;
        RECT 2898.070 2429.000 2898.390 2429.060 ;
      LAYER via ;
        RECT 1984.540 2429.000 1984.800 2429.260 ;
        RECT 2898.100 2429.000 2898.360 2429.260 ;
      LAYER met2 ;
        RECT 2898.090 2433.875 2898.370 2434.245 ;
        RECT 2898.160 2429.290 2898.300 2433.875 ;
        RECT 1984.540 2428.970 1984.800 2429.290 ;
        RECT 2898.100 2428.970 2898.360 2429.290 ;
        RECT 1984.600 1064.045 1984.740 2428.970 ;
        RECT 1984.530 1063.675 1984.810 1064.045 ;
      LAYER via2 ;
        RECT 2898.090 2433.920 2898.370 2434.200 ;
        RECT 1984.530 1063.720 1984.810 1064.000 ;
      LAYER met3 ;
        RECT 2898.065 2434.210 2898.395 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2898.065 2433.910 2924.800 2434.210 ;
        RECT 2898.065 2433.895 2898.395 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
        RECT 1966.720 1064.010 1970.720 1064.200 ;
        RECT 1984.505 1064.010 1984.835 1064.025 ;
        RECT 1966.720 1063.710 1984.835 1064.010 ;
        RECT 1966.720 1063.600 1970.720 1063.710 ;
        RECT 1984.505 1063.695 1984.835 1063.710 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1759.110 2663.800 1759.430 2663.860 ;
        RECT 2900.830 2663.800 2901.150 2663.860 ;
        RECT 1759.110 2663.660 2901.150 2663.800 ;
        RECT 1759.110 2663.600 1759.430 2663.660 ;
        RECT 2900.830 2663.600 2901.150 2663.660 ;
      LAYER via ;
        RECT 1759.140 2663.600 1759.400 2663.860 ;
        RECT 2900.860 2663.600 2901.120 2663.860 ;
      LAYER met2 ;
        RECT 2900.850 2669.155 2901.130 2669.525 ;
        RECT 2900.920 2663.890 2901.060 2669.155 ;
        RECT 1759.140 2663.570 1759.400 2663.890 ;
        RECT 2900.860 2663.570 2901.120 2663.890 ;
        RECT 1759.200 951.165 1759.340 2663.570 ;
        RECT 1759.130 950.795 1759.410 951.165 ;
      LAYER via2 ;
        RECT 2900.850 2669.200 2901.130 2669.480 ;
        RECT 1759.130 950.840 1759.410 951.120 ;
      LAYER met3 ;
        RECT 2900.825 2669.490 2901.155 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2900.825 2669.190 2924.800 2669.490 ;
        RECT 2900.825 2669.175 2901.155 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
        RECT 1759.105 951.130 1759.435 951.145 ;
        RECT 1770.720 951.130 1774.720 951.320 ;
        RECT 1759.105 950.830 1774.720 951.130 ;
        RECT 1759.105 950.815 1759.435 950.830 ;
        RECT 1770.720 950.720 1774.720 950.830 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1984.050 2898.400 1984.370 2898.460 ;
        RECT 2900.830 2898.400 2901.150 2898.460 ;
        RECT 1984.050 2898.260 2901.150 2898.400 ;
        RECT 1984.050 2898.200 1984.370 2898.260 ;
        RECT 2900.830 2898.200 2901.150 2898.260 ;
      LAYER via ;
        RECT 1984.080 2898.200 1984.340 2898.460 ;
        RECT 2900.860 2898.200 2901.120 2898.460 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2898.490 2901.060 2903.755 ;
        RECT 1984.080 2898.170 1984.340 2898.490 ;
        RECT 2900.860 2898.170 2901.120 2898.490 ;
        RECT 1984.140 959.325 1984.280 2898.170 ;
        RECT 1984.070 958.955 1984.350 959.325 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
        RECT 1984.070 959.000 1984.350 959.280 ;
      LAYER met3 ;
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
        RECT 1966.720 959.290 1970.720 959.480 ;
        RECT 1984.045 959.290 1984.375 959.305 ;
        RECT 1966.720 958.990 1984.375 959.290 ;
        RECT 1966.720 958.880 1970.720 958.990 ;
        RECT 1984.045 958.975 1984.375 958.990 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1959.210 3133.000 1959.530 3133.060 ;
        RECT 2900.830 3133.000 2901.150 3133.060 ;
        RECT 1959.210 3132.860 2901.150 3133.000 ;
        RECT 1959.210 3132.800 1959.530 3132.860 ;
        RECT 2900.830 3132.800 2901.150 3132.860 ;
      LAYER via ;
        RECT 1959.240 3132.800 1959.500 3133.060 ;
        RECT 2900.860 3132.800 2901.120 3133.060 ;
      LAYER met2 ;
        RECT 2900.850 3138.355 2901.130 3138.725 ;
        RECT 2900.920 3133.090 2901.060 3138.355 ;
        RECT 1959.240 3132.770 1959.500 3133.090 ;
        RECT 2900.860 3132.770 2901.120 3133.090 ;
        RECT 1956.550 1119.010 1956.830 1120.000 ;
        RECT 1959.300 1119.010 1959.440 3132.770 ;
        RECT 1956.550 1118.870 1959.440 1119.010 ;
        RECT 1956.550 1116.000 1956.830 1118.870 ;
      LAYER via2 ;
        RECT 2900.850 3138.400 2901.130 3138.680 ;
      LAYER met3 ;
        RECT 2900.825 3138.690 2901.155 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.825 3138.390 2924.800 3138.690 ;
        RECT 2900.825 3138.375 2901.155 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1983.590 3367.600 1983.910 3367.660 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 1983.590 3367.460 2901.150 3367.600 ;
        RECT 1983.590 3367.400 1983.910 3367.460 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
      LAYER via ;
        RECT 1983.620 3367.400 1983.880 3367.660 ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 1983.620 3367.370 1983.880 3367.690 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
        RECT 1983.680 1030.045 1983.820 3367.370 ;
        RECT 1983.610 1029.675 1983.890 1030.045 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
        RECT 1983.610 1029.720 1983.890 1030.000 ;
      LAYER met3 ;
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
        RECT 1966.720 1030.010 1970.720 1030.200 ;
        RECT 1983.585 1030.010 1983.915 1030.025 ;
        RECT 1966.720 1029.710 1983.915 1030.010 ;
        RECT 1966.720 1029.600 1970.720 1029.710 ;
        RECT 1983.585 1029.695 1983.915 1029.710 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1855.710 3501.560 1856.030 3501.620 ;
        RECT 2798.250 3501.560 2798.570 3501.620 ;
        RECT 1855.710 3501.420 2798.570 3501.560 ;
        RECT 1855.710 3501.360 1856.030 3501.420 ;
        RECT 2798.250 3501.360 2798.570 3501.420 ;
        RECT 1849.730 1132.100 1850.050 1132.160 ;
        RECT 1855.710 1132.100 1856.030 1132.160 ;
        RECT 1849.730 1131.960 1856.030 1132.100 ;
        RECT 1849.730 1131.900 1850.050 1131.960 ;
        RECT 1855.710 1131.900 1856.030 1131.960 ;
      LAYER via ;
        RECT 1855.740 3501.360 1856.000 3501.620 ;
        RECT 2798.280 3501.360 2798.540 3501.620 ;
        RECT 1849.760 1131.900 1850.020 1132.160 ;
        RECT 1855.740 1131.900 1856.000 1132.160 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3501.650 2798.480 3517.600 ;
        RECT 1855.740 3501.330 1856.000 3501.650 ;
        RECT 2798.280 3501.330 2798.540 3501.650 ;
        RECT 1855.800 1132.190 1855.940 3501.330 ;
        RECT 1849.760 1131.870 1850.020 1132.190 ;
        RECT 1855.740 1131.870 1856.000 1132.190 ;
        RECT 1849.820 1120.000 1849.960 1131.870 ;
        RECT 1849.820 1119.620 1850.110 1120.000 ;
        RECT 1849.830 1116.000 1850.110 1119.620 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1938.510 3501.900 1938.830 3501.960 ;
        RECT 2473.950 3501.900 2474.270 3501.960 ;
        RECT 1938.510 3501.760 2474.270 3501.900 ;
        RECT 1938.510 3501.700 1938.830 3501.760 ;
        RECT 2473.950 3501.700 2474.270 3501.760 ;
        RECT 1932.530 1132.100 1932.850 1132.160 ;
        RECT 1938.510 1132.100 1938.830 1132.160 ;
        RECT 1932.530 1131.960 1938.830 1132.100 ;
        RECT 1932.530 1131.900 1932.850 1131.960 ;
        RECT 1938.510 1131.900 1938.830 1131.960 ;
      LAYER via ;
        RECT 1938.540 3501.700 1938.800 3501.960 ;
        RECT 2473.980 3501.700 2474.240 3501.960 ;
        RECT 1932.560 1131.900 1932.820 1132.160 ;
        RECT 1938.540 1131.900 1938.800 1132.160 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3501.990 2474.180 3517.600 ;
        RECT 1938.540 3501.670 1938.800 3501.990 ;
        RECT 2473.980 3501.670 2474.240 3501.990 ;
        RECT 1938.600 1132.190 1938.740 3501.670 ;
        RECT 1932.560 1131.870 1932.820 1132.190 ;
        RECT 1938.540 1131.870 1938.800 1132.190 ;
        RECT 1932.620 1120.000 1932.760 1131.870 ;
        RECT 1932.620 1119.620 1932.910 1120.000 ;
        RECT 1932.630 1116.000 1932.910 1119.620 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1890.210 3502.240 1890.530 3502.300 ;
        RECT 2149.190 3502.240 2149.510 3502.300 ;
        RECT 1890.210 3502.100 2149.510 3502.240 ;
        RECT 1890.210 3502.040 1890.530 3502.100 ;
        RECT 2149.190 3502.040 2149.510 3502.100 ;
        RECT 1885.610 1132.100 1885.930 1132.160 ;
        RECT 1890.210 1132.100 1890.530 1132.160 ;
        RECT 1885.610 1131.960 1890.530 1132.100 ;
        RECT 1885.610 1131.900 1885.930 1131.960 ;
        RECT 1890.210 1131.900 1890.530 1131.960 ;
      LAYER via ;
        RECT 1890.240 3502.040 1890.500 3502.300 ;
        RECT 2149.220 3502.040 2149.480 3502.300 ;
        RECT 1885.640 1131.900 1885.900 1132.160 ;
        RECT 1890.240 1131.900 1890.500 1132.160 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3502.330 2149.420 3517.600 ;
        RECT 1890.240 3502.010 1890.500 3502.330 ;
        RECT 2149.220 3502.010 2149.480 3502.330 ;
        RECT 1890.300 1132.190 1890.440 3502.010 ;
        RECT 1885.640 1131.870 1885.900 1132.190 ;
        RECT 1890.240 1131.870 1890.500 1132.190 ;
        RECT 1885.700 1120.000 1885.840 1131.870 ;
        RECT 1885.700 1119.620 1885.990 1120.000 ;
        RECT 1885.710 1116.000 1885.990 1119.620 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1773.830 3501.560 1774.150 3501.620 ;
        RECT 1824.890 3501.560 1825.210 3501.620 ;
        RECT 1773.830 3501.420 1825.210 3501.560 ;
        RECT 1773.830 3501.360 1774.150 3501.420 ;
        RECT 1824.890 3501.360 1825.210 3501.420 ;
      LAYER via ;
        RECT 1773.860 3501.360 1774.120 3501.620 ;
        RECT 1824.920 3501.360 1825.180 3501.620 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3501.650 1825.120 3517.600 ;
        RECT 1773.860 3501.330 1774.120 3501.650 ;
        RECT 1824.920 3501.330 1825.180 3501.650 ;
        RECT 1773.920 924.530 1774.060 3501.330 ;
        RECT 1773.920 924.390 1778.660 924.530 ;
        RECT 1778.520 923.850 1778.660 924.390 ;
        RECT 1779.910 923.850 1780.190 924.000 ;
        RECT 1778.520 923.710 1780.190 923.850 ;
        RECT 1779.910 920.000 1780.190 923.710 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1775.745 906.185 1775.915 908.735 ;
      LAYER mcon ;
        RECT 1775.745 908.565 1775.915 908.735 ;
      LAYER met1 ;
        RECT 1500.590 3498.500 1500.910 3498.560 ;
        RECT 1503.810 3498.500 1504.130 3498.560 ;
        RECT 1500.590 3498.360 1504.130 3498.500 ;
        RECT 1500.590 3498.300 1500.910 3498.360 ;
        RECT 1503.810 3498.300 1504.130 3498.360 ;
        RECT 1503.810 908.720 1504.130 908.780 ;
        RECT 1775.685 908.720 1775.975 908.765 ;
        RECT 1503.810 908.580 1775.975 908.720 ;
        RECT 1503.810 908.520 1504.130 908.580 ;
        RECT 1775.685 908.535 1775.975 908.580 ;
        RECT 1775.685 906.340 1775.975 906.385 ;
        RECT 1814.770 906.340 1815.090 906.400 ;
        RECT 1775.685 906.200 1815.090 906.340 ;
        RECT 1775.685 906.155 1775.975 906.200 ;
        RECT 1814.770 906.140 1815.090 906.200 ;
      LAYER via ;
        RECT 1500.620 3498.300 1500.880 3498.560 ;
        RECT 1503.840 3498.300 1504.100 3498.560 ;
        RECT 1503.840 908.520 1504.100 908.780 ;
        RECT 1814.800 906.140 1815.060 906.400 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3498.590 1500.820 3517.600 ;
        RECT 1500.620 3498.270 1500.880 3498.590 ;
        RECT 1503.840 3498.270 1504.100 3498.590 ;
        RECT 1503.900 908.810 1504.040 3498.270 ;
        RECT 1814.870 920.380 1815.150 924.000 ;
        RECT 1814.860 920.000 1815.150 920.380 ;
        RECT 1503.840 908.490 1504.100 908.810 ;
        RECT 1814.860 906.430 1815.000 920.000 ;
        RECT 1814.800 906.110 1815.060 906.430 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 322.060 2924.800 323.260 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3410.620 2.400 3411.820 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3123.660 2.400 3124.860 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2836.020 2.400 2837.220 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2549.060 2.400 2550.260 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2261.420 2.400 2262.620 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1974.460 2.400 1975.660 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 556.660 2924.800 557.860 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1686.820 2.400 1688.020 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1471.260 2.400 1472.460 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1255.700 2.400 1256.900 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1040.140 2.400 1041.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 824.580 2.400 825.780 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 609.700 2.400 610.900 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 394.140 2.400 395.340 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 178.580 2.400 179.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 791.260 2924.800 792.460 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1025.860 2924.800 1027.060 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1260.460 2924.800 1261.660 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1495.060 2924.800 1496.260 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1729.660 2924.800 1730.860 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1758.650 1960.000 1758.970 1960.060 ;
        RECT 2899.450 1960.000 2899.770 1960.060 ;
        RECT 1758.650 1959.860 2899.770 1960.000 ;
        RECT 1758.650 1959.800 1758.970 1959.860 ;
        RECT 2899.450 1959.800 2899.770 1959.860 ;
      LAYER via ;
        RECT 1758.680 1959.800 1758.940 1960.060 ;
        RECT 2899.480 1959.800 2899.740 1960.060 ;
      LAYER met2 ;
        RECT 2899.470 1964.675 2899.750 1965.045 ;
        RECT 2899.540 1960.090 2899.680 1964.675 ;
        RECT 1758.680 1959.770 1758.940 1960.090 ;
        RECT 2899.480 1959.770 2899.740 1960.090 ;
        RECT 1758.740 1072.205 1758.880 1959.770 ;
        RECT 1758.670 1071.835 1758.950 1072.205 ;
      LAYER via2 ;
        RECT 2899.470 1964.720 2899.750 1965.000 ;
        RECT 1758.670 1071.880 1758.950 1072.160 ;
      LAYER met3 ;
        RECT 2899.445 1965.010 2899.775 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2899.445 1964.710 2924.800 1965.010 ;
        RECT 2899.445 1964.695 2899.775 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
        RECT 1758.645 1072.170 1758.975 1072.185 ;
        RECT 1770.720 1072.170 1774.720 1072.360 ;
        RECT 1758.645 1071.870 1774.720 1072.170 ;
        RECT 1758.645 1071.855 1758.975 1071.870 ;
        RECT 1770.720 1071.760 1774.720 1071.870 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1976.690 2194.600 1977.010 2194.660 ;
        RECT 2898.070 2194.600 2898.390 2194.660 ;
        RECT 1976.690 2194.460 2898.390 2194.600 ;
        RECT 1976.690 2194.400 1977.010 2194.460 ;
        RECT 2898.070 2194.400 2898.390 2194.460 ;
        RECT 1826.730 909.060 1827.050 909.120 ;
        RECT 1976.690 909.060 1977.010 909.120 ;
        RECT 1826.730 908.920 1977.010 909.060 ;
        RECT 1826.730 908.860 1827.050 908.920 ;
        RECT 1976.690 908.860 1977.010 908.920 ;
      LAYER via ;
        RECT 1976.720 2194.400 1976.980 2194.660 ;
        RECT 2898.100 2194.400 2898.360 2194.660 ;
        RECT 1826.760 908.860 1827.020 909.120 ;
        RECT 1976.720 908.860 1976.980 909.120 ;
      LAYER met2 ;
        RECT 2898.090 2199.275 2898.370 2199.645 ;
        RECT 2898.160 2194.690 2898.300 2199.275 ;
        RECT 1976.720 2194.370 1976.980 2194.690 ;
        RECT 2898.100 2194.370 2898.360 2194.690 ;
        RECT 1826.830 920.380 1827.110 924.000 ;
        RECT 1826.820 920.000 1827.110 920.380 ;
        RECT 1826.820 909.150 1826.960 920.000 ;
        RECT 1976.780 909.150 1976.920 2194.370 ;
        RECT 1826.760 908.830 1827.020 909.150 ;
        RECT 1976.720 908.830 1976.980 909.150 ;
      LAYER via2 ;
        RECT 2898.090 2199.320 2898.370 2199.600 ;
      LAYER met3 ;
        RECT 2898.065 2199.610 2898.395 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2898.065 2199.310 2924.800 2199.610 ;
        RECT 2898.065 2199.295 2898.395 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 204.420 2924.800 205.620 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 439.020 2924.800 440.220 ;
    END
  END io_oeb[1]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1830.300 2.400 1831.500 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 673.620 2924.800 674.820 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1543.340 2.400 1544.540 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1327.780 2.400 1328.980 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1112.220 2.400 1113.420 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 896.660 2.400 897.860 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 681.100 2.400 682.300 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 465.540 2.400 466.740 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 249.980 2.400 251.180 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 35.100 2.400 36.300 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 908.900 2924.800 910.100 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1143.500 2924.800 1144.700 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1378.100 2924.800 1379.300 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1612.700 2924.800 1613.900 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1847.300 2924.800 1848.500 ;
    END
  END io_oeb[7]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 145.940 2924.800 147.140 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2492.620 2924.800 2493.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2727.220 2924.800 2728.420 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2961.820 2924.800 2963.020 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3196.420 2924.800 3197.620 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3431.020 2924.800 3432.220 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 380.540 2924.800 381.740 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1094.870 3502.580 1095.190 3502.640 ;
        RECT 1762.790 3502.580 1763.110 3502.640 ;
        RECT 1094.870 3502.440 1763.110 3502.580 ;
        RECT 1094.870 3502.380 1095.190 3502.440 ;
        RECT 1762.790 3502.380 1763.110 3502.440 ;
        RECT 1762.790 907.700 1763.110 907.760 ;
        RECT 1897.570 907.700 1897.890 907.760 ;
        RECT 1762.790 907.560 1897.890 907.700 ;
        RECT 1762.790 907.500 1763.110 907.560 ;
        RECT 1897.570 907.500 1897.890 907.560 ;
      LAYER via ;
        RECT 1094.900 3502.380 1095.160 3502.640 ;
        RECT 1762.820 3502.380 1763.080 3502.640 ;
        RECT 1762.820 907.500 1763.080 907.760 ;
        RECT 1897.600 907.500 1897.860 907.760 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3502.670 1095.100 3517.600 ;
        RECT 1094.900 3502.350 1095.160 3502.670 ;
        RECT 1762.820 3502.350 1763.080 3502.670 ;
        RECT 1762.880 907.790 1763.020 3502.350 ;
        RECT 1897.670 920.380 1897.950 924.000 ;
        RECT 1897.660 920.000 1897.950 920.380 ;
        RECT 1897.660 907.790 1897.800 920.000 ;
        RECT 1762.820 907.470 1763.080 907.790 ;
        RECT 1897.600 907.470 1897.860 907.790 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 770.570 3502.240 770.890 3502.300 ;
        RECT 1493.690 3502.240 1494.010 3502.300 ;
        RECT 770.570 3502.100 1494.010 3502.240 ;
        RECT 770.570 3502.040 770.890 3502.100 ;
        RECT 1493.690 3502.040 1494.010 3502.100 ;
        RECT 1493.690 1041.660 1494.010 1041.720 ;
        RECT 1752.670 1041.660 1752.990 1041.720 ;
        RECT 1493.690 1041.520 1752.990 1041.660 ;
        RECT 1493.690 1041.460 1494.010 1041.520 ;
        RECT 1752.670 1041.460 1752.990 1041.520 ;
      LAYER via ;
        RECT 770.600 3502.040 770.860 3502.300 ;
        RECT 1493.720 3502.040 1493.980 3502.300 ;
        RECT 1493.720 1041.460 1493.980 1041.720 ;
        RECT 1752.700 1041.460 1752.960 1041.720 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3502.330 770.800 3517.600 ;
        RECT 770.600 3502.010 770.860 3502.330 ;
        RECT 1493.720 3502.010 1493.980 3502.330 ;
        RECT 1493.780 1041.750 1493.920 3502.010 ;
        RECT 1493.720 1041.430 1493.980 1041.750 ;
        RECT 1752.700 1041.430 1752.960 1041.750 ;
        RECT 1752.760 1038.205 1752.900 1041.430 ;
        RECT 1752.690 1037.835 1752.970 1038.205 ;
      LAYER via2 ;
        RECT 1752.690 1037.880 1752.970 1038.160 ;
      LAYER met3 ;
        RECT 1752.665 1038.170 1752.995 1038.185 ;
        RECT 1770.720 1038.170 1774.720 1038.360 ;
        RECT 1752.665 1037.870 1774.720 1038.170 ;
        RECT 1752.665 1037.855 1752.995 1037.870 ;
        RECT 1770.720 1037.760 1774.720 1037.870 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3501.900 446.130 3501.960 ;
        RECT 1783.490 3501.900 1783.810 3501.960 ;
        RECT 445.810 3501.760 1783.810 3501.900 ;
        RECT 445.810 3501.700 446.130 3501.760 ;
        RECT 1783.490 3501.700 1783.810 3501.760 ;
        RECT 1783.490 1135.500 1783.810 1135.560 ;
        RECT 1873.650 1135.500 1873.970 1135.560 ;
        RECT 1783.490 1135.360 1873.970 1135.500 ;
        RECT 1783.490 1135.300 1783.810 1135.360 ;
        RECT 1873.650 1135.300 1873.970 1135.360 ;
      LAYER via ;
        RECT 445.840 3501.700 446.100 3501.960 ;
        RECT 1783.520 3501.700 1783.780 3501.960 ;
        RECT 1783.520 1135.300 1783.780 1135.560 ;
        RECT 1873.680 1135.300 1873.940 1135.560 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3501.990 446.040 3517.600 ;
        RECT 445.840 3501.670 446.100 3501.990 ;
        RECT 1783.520 3501.670 1783.780 3501.990 ;
        RECT 1783.580 1135.590 1783.720 3501.670 ;
        RECT 1783.520 1135.270 1783.780 1135.590 ;
        RECT 1873.680 1135.270 1873.940 1135.590 ;
        RECT 1873.740 1120.000 1873.880 1135.270 ;
        RECT 1873.740 1119.620 1874.030 1120.000 ;
        RECT 1873.750 1116.000 1874.030 1119.620 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3501.560 121.830 3501.620 ;
        RECT 1507.490 3501.560 1507.810 3501.620 ;
        RECT 121.510 3501.420 1507.810 3501.560 ;
        RECT 121.510 3501.360 121.830 3501.420 ;
        RECT 1507.490 3501.360 1507.810 3501.420 ;
        RECT 1507.490 972.640 1507.810 972.700 ;
        RECT 1752.670 972.640 1752.990 972.700 ;
        RECT 1507.490 972.500 1752.990 972.640 ;
        RECT 1507.490 972.440 1507.810 972.500 ;
        RECT 1752.670 972.440 1752.990 972.500 ;
      LAYER via ;
        RECT 121.540 3501.360 121.800 3501.620 ;
        RECT 1507.520 3501.360 1507.780 3501.620 ;
        RECT 1507.520 972.440 1507.780 972.700 ;
        RECT 1752.700 972.440 1752.960 972.700 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3501.650 121.740 3517.600 ;
        RECT 121.540 3501.330 121.800 3501.650 ;
        RECT 1507.520 3501.330 1507.780 3501.650 ;
        RECT 1507.580 972.730 1507.720 3501.330 ;
        RECT 1507.520 972.410 1507.780 972.730 ;
        RECT 1752.700 972.410 1752.960 972.730 ;
        RECT 1752.760 967.485 1752.900 972.410 ;
        RECT 1752.690 967.115 1752.970 967.485 ;
      LAYER via2 ;
        RECT 1752.690 967.160 1752.970 967.440 ;
      LAYER met3 ;
        RECT 1752.665 967.450 1752.995 967.465 ;
        RECT 1770.720 967.450 1774.720 967.640 ;
        RECT 1752.665 967.150 1774.720 967.450 ;
        RECT 1752.665 967.135 1752.995 967.150 ;
        RECT 1770.720 967.040 1774.720 967.150 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3339.720 17.410 3339.780 ;
        RECT 1514.390 3339.720 1514.710 3339.780 ;
        RECT 17.090 3339.580 1514.710 3339.720 ;
        RECT 17.090 3339.520 17.410 3339.580 ;
        RECT 1514.390 3339.520 1514.710 3339.580 ;
        RECT 1514.390 931.500 1514.710 931.560 ;
        RECT 1968.870 931.500 1969.190 931.560 ;
        RECT 1514.390 931.360 1969.190 931.500 ;
        RECT 1514.390 931.300 1514.710 931.360 ;
        RECT 1968.870 931.300 1969.190 931.360 ;
      LAYER via ;
        RECT 17.120 3339.520 17.380 3339.780 ;
        RECT 1514.420 3339.520 1514.680 3339.780 ;
        RECT 1514.420 931.300 1514.680 931.560 ;
        RECT 1968.900 931.300 1969.160 931.560 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.120 3339.490 17.380 3339.635 ;
        RECT 1514.420 3339.490 1514.680 3339.810 ;
        RECT 1514.480 931.590 1514.620 3339.490 ;
        RECT 1514.420 931.270 1514.680 931.590 ;
        RECT 1968.900 931.270 1969.160 931.590 ;
        RECT 1968.960 928.045 1969.100 931.270 ;
        RECT 1968.890 927.675 1969.170 928.045 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
        RECT 1968.890 927.720 1969.170 928.000 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
        RECT 1968.865 928.010 1969.195 928.025 ;
        RECT 1968.865 927.695 1969.410 928.010 ;
        RECT 1969.110 925.480 1969.410 927.695 ;
        RECT 1966.720 924.880 1970.720 925.480 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3050.040 17.410 3050.100 ;
        RECT 1967.950 3050.040 1968.270 3050.100 ;
        RECT 17.090 3049.900 1968.270 3050.040 ;
        RECT 17.090 3049.840 17.410 3049.900 ;
        RECT 1967.950 3049.840 1968.270 3049.900 ;
      LAYER via ;
        RECT 17.120 3049.840 17.380 3050.100 ;
        RECT 1967.980 3049.840 1968.240 3050.100 ;
      LAYER met2 ;
        RECT 17.110 3051.995 17.390 3052.365 ;
        RECT 17.180 3050.130 17.320 3051.995 ;
        RECT 17.120 3049.810 17.380 3050.130 ;
        RECT 1967.980 3049.810 1968.240 3050.130 ;
        RECT 1968.040 1013.610 1968.180 3049.810 ;
        RECT 1968.430 1013.610 1968.710 1013.725 ;
        RECT 1968.040 1013.470 1968.710 1013.610 ;
        RECT 1968.430 1013.355 1968.710 1013.470 ;
      LAYER via2 ;
        RECT 17.110 3052.040 17.390 3052.320 ;
        RECT 1968.430 1013.400 1968.710 1013.680 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 17.085 3052.330 17.415 3052.345 ;
        RECT -4.800 3052.030 17.415 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 17.085 3052.015 17.415 3052.030 ;
        RECT 1968.405 1013.690 1968.735 1013.705 ;
        RECT 1968.190 1013.375 1968.735 1013.690 ;
        RECT 1968.190 1012.520 1968.490 1013.375 ;
        RECT 1966.720 1011.920 1970.720 1012.520 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2760.360 16.030 2760.420 ;
        RECT 1797.290 2760.360 1797.610 2760.420 ;
        RECT 15.710 2760.220 1797.610 2760.360 ;
        RECT 15.710 2760.160 16.030 2760.220 ;
        RECT 1797.290 2760.160 1797.610 2760.220 ;
        RECT 1797.290 1132.100 1797.610 1132.160 ;
        RECT 1814.770 1132.100 1815.090 1132.160 ;
        RECT 1797.290 1131.960 1815.090 1132.100 ;
        RECT 1797.290 1131.900 1797.610 1131.960 ;
        RECT 1814.770 1131.900 1815.090 1131.960 ;
      LAYER via ;
        RECT 15.740 2760.160 16.000 2760.420 ;
        RECT 1797.320 2760.160 1797.580 2760.420 ;
        RECT 1797.320 1131.900 1797.580 1132.160 ;
        RECT 1814.800 1131.900 1815.060 1132.160 ;
      LAYER met2 ;
        RECT 15.730 2765.035 16.010 2765.405 ;
        RECT 15.800 2760.450 15.940 2765.035 ;
        RECT 15.740 2760.130 16.000 2760.450 ;
        RECT 1797.320 2760.130 1797.580 2760.450 ;
        RECT 1797.380 1132.190 1797.520 2760.130 ;
        RECT 1797.320 1131.870 1797.580 1132.190 ;
        RECT 1814.800 1131.870 1815.060 1132.190 ;
        RECT 1814.860 1120.000 1815.000 1131.870 ;
        RECT 1814.860 1119.620 1815.150 1120.000 ;
        RECT 1814.870 1116.000 1815.150 1119.620 ;
      LAYER via2 ;
        RECT 15.730 2765.080 16.010 2765.360 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 15.705 2765.370 16.035 2765.385 ;
        RECT -4.800 2765.070 16.035 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 15.705 2765.055 16.035 2765.070 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2477.480 17.410 2477.540 ;
        RECT 1521.290 2477.480 1521.610 2477.540 ;
        RECT 17.090 2477.340 1521.610 2477.480 ;
        RECT 17.090 2477.280 17.410 2477.340 ;
        RECT 1521.290 2477.280 1521.610 2477.340 ;
        RECT 1521.290 1135.160 1521.610 1135.220 ;
        RECT 1802.810 1135.160 1803.130 1135.220 ;
        RECT 1521.290 1135.020 1803.130 1135.160 ;
        RECT 1521.290 1134.960 1521.610 1135.020 ;
        RECT 1802.810 1134.960 1803.130 1135.020 ;
      LAYER via ;
        RECT 17.120 2477.280 17.380 2477.540 ;
        RECT 1521.320 2477.280 1521.580 2477.540 ;
        RECT 1521.320 1134.960 1521.580 1135.220 ;
        RECT 1802.840 1134.960 1803.100 1135.220 ;
      LAYER met2 ;
        RECT 17.110 2477.395 17.390 2477.765 ;
        RECT 17.120 2477.250 17.380 2477.395 ;
        RECT 1521.320 2477.250 1521.580 2477.570 ;
        RECT 1521.380 1135.250 1521.520 2477.250 ;
        RECT 1521.320 1134.930 1521.580 1135.250 ;
        RECT 1802.840 1134.930 1803.100 1135.250 ;
        RECT 1802.900 1120.000 1803.040 1134.930 ;
        RECT 1802.900 1119.620 1803.190 1120.000 ;
        RECT 1802.910 1116.000 1803.190 1119.620 ;
      LAYER via2 ;
        RECT 17.110 2477.440 17.390 2477.720 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 17.085 2477.730 17.415 2477.745 ;
        RECT -4.800 2477.430 17.415 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 17.085 2477.415 17.415 2477.430 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2187.460 17.870 2187.520 ;
        RECT 1528.190 2187.460 1528.510 2187.520 ;
        RECT 17.550 2187.320 1528.510 2187.460 ;
        RECT 17.550 2187.260 17.870 2187.320 ;
        RECT 1528.190 2187.260 1528.510 2187.320 ;
        RECT 1528.190 1007.320 1528.510 1007.380 ;
        RECT 1752.670 1007.320 1752.990 1007.380 ;
        RECT 1528.190 1007.180 1752.990 1007.320 ;
        RECT 1528.190 1007.120 1528.510 1007.180 ;
        RECT 1752.670 1007.120 1752.990 1007.180 ;
      LAYER via ;
        RECT 17.580 2187.260 17.840 2187.520 ;
        RECT 1528.220 2187.260 1528.480 2187.520 ;
        RECT 1528.220 1007.120 1528.480 1007.380 ;
        RECT 1752.700 1007.120 1752.960 1007.380 ;
      LAYER met2 ;
        RECT 17.570 2189.755 17.850 2190.125 ;
        RECT 17.640 2187.550 17.780 2189.755 ;
        RECT 17.580 2187.230 17.840 2187.550 ;
        RECT 1528.220 2187.230 1528.480 2187.550 ;
        RECT 1528.280 1007.410 1528.420 2187.230 ;
        RECT 1528.220 1007.090 1528.480 1007.410 ;
        RECT 1752.700 1007.090 1752.960 1007.410 ;
        RECT 1752.760 1002.845 1752.900 1007.090 ;
        RECT 1752.690 1002.475 1752.970 1002.845 ;
      LAYER via2 ;
        RECT 17.570 2189.800 17.850 2190.080 ;
        RECT 1752.690 1002.520 1752.970 1002.800 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 17.545 2190.090 17.875 2190.105 ;
        RECT -4.800 2189.790 17.875 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 17.545 2189.775 17.875 2189.790 ;
        RECT 1752.665 1002.810 1752.995 1002.825 ;
        RECT 1770.720 1002.810 1774.720 1003.000 ;
        RECT 1752.665 1002.510 1774.720 1002.810 ;
        RECT 1752.665 1002.495 1752.995 1002.510 ;
        RECT 1770.720 1002.400 1774.720 1002.510 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1902.380 2.400 1903.580 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 615.140 2924.800 616.340 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1614.740 2.400 1615.940 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1184.300 2.400 1185.500 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 968.740 2.400 969.940 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 753.180 2.400 754.380 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 537.620 2.400 538.820 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 322.060 2.400 323.260 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 106.500 2.400 107.700 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 849.740 2924.800 850.940 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1084.340 2924.800 1085.540 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1318.940 2924.800 1320.140 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1553.540 2924.800 1554.740 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1788.820 2924.800 1790.020 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2023.420 2924.800 2024.620 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2258.020 2924.800 2259.220 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 3504.960 1338.530 3505.020 ;
        RECT 1662.510 3504.960 1662.830 3505.020 ;
        RECT 1987.270 3504.960 1987.590 3505.020 ;
        RECT 2311.570 3504.960 2311.890 3505.020 ;
        RECT 2635.870 3504.960 2636.190 3505.020 ;
        RECT 1338.210 3504.820 2636.190 3504.960 ;
        RECT 1338.210 3504.760 1338.530 3504.820 ;
        RECT 1662.510 3504.760 1662.830 3504.820 ;
        RECT 1987.270 3504.760 1987.590 3504.820 ;
        RECT 2311.570 3504.760 2311.890 3504.820 ;
        RECT 2635.870 3504.760 2636.190 3504.820 ;
        RECT 2635.870 3501.900 2636.190 3501.960 ;
        RECT 2902.210 3501.900 2902.530 3501.960 ;
        RECT 2635.870 3501.760 2902.530 3501.900 ;
        RECT 2635.870 3501.700 2636.190 3501.760 ;
        RECT 2902.210 3501.700 2902.530 3501.760 ;
        RECT 1986.810 1048.800 1987.130 1048.860 ;
        RECT 2901.290 1048.800 2901.610 1048.860 ;
        RECT 1986.810 1048.660 2901.610 1048.800 ;
        RECT 1986.810 1048.600 1987.130 1048.660 ;
        RECT 2901.290 1048.600 2901.610 1048.660 ;
      LAYER via ;
        RECT 1338.240 3504.760 1338.500 3505.020 ;
        RECT 1662.540 3504.760 1662.800 3505.020 ;
        RECT 1987.300 3504.760 1987.560 3505.020 ;
        RECT 2311.600 3504.760 2311.860 3505.020 ;
        RECT 2635.900 3504.760 2636.160 3505.020 ;
        RECT 2635.900 3501.700 2636.160 3501.960 ;
        RECT 2902.240 3501.700 2902.500 3501.960 ;
        RECT 1986.840 1048.600 1987.100 1048.860 ;
        RECT 2901.320 1048.600 2901.580 1048.860 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 1338.300 3505.050 1338.440 3517.600 ;
        RECT 1662.600 3505.050 1662.740 3517.600 ;
        RECT 1987.360 3505.050 1987.500 3517.600 ;
        RECT 2311.660 3505.050 2311.800 3517.600 ;
        RECT 2635.960 3505.050 2636.100 3517.600 ;
        RECT 1338.240 3504.730 1338.500 3505.050 ;
        RECT 1662.540 3504.730 1662.800 3505.050 ;
        RECT 1987.300 3504.730 1987.560 3505.050 ;
        RECT 2311.600 3504.730 2311.860 3505.050 ;
        RECT 2635.900 3504.730 2636.160 3505.050 ;
        RECT 2635.960 3501.990 2636.100 3504.730 ;
        RECT 2635.900 3501.670 2636.160 3501.990 ;
        RECT 2902.240 3501.670 2902.500 3501.990 ;
        RECT 2902.300 3490.285 2902.440 3501.670 ;
        RECT 2902.230 3489.915 2902.510 3490.285 ;
        RECT 2904.530 3489.915 2904.810 3490.285 ;
        RECT 2904.600 3255.685 2904.740 3489.915 ;
        RECT 2904.530 3255.315 2904.810 3255.685 ;
        RECT 2904.600 3021.085 2904.740 3255.315 ;
        RECT 2904.530 3020.715 2904.810 3021.085 ;
        RECT 2904.600 2786.485 2904.740 3020.715 ;
        RECT 2904.530 2786.115 2904.810 2786.485 ;
        RECT 2904.600 2551.885 2904.740 2786.115 ;
        RECT 2904.530 2551.515 2904.810 2551.885 ;
        RECT 2904.600 2317.285 2904.740 2551.515 ;
        RECT 2904.530 2316.915 2904.810 2317.285 ;
        RECT 2904.600 2082.685 2904.740 2316.915 ;
        RECT 2901.310 2082.315 2901.590 2082.685 ;
        RECT 2904.530 2082.315 2904.810 2082.685 ;
        RECT 2901.380 1048.890 2901.520 2082.315 ;
        RECT 1986.840 1048.570 1987.100 1048.890 ;
        RECT 2901.320 1048.570 2901.580 1048.890 ;
        RECT 1986.900 1046.365 1987.040 1048.570 ;
        RECT 1986.830 1045.995 1987.110 1046.365 ;
      LAYER via2 ;
        RECT 2902.230 3489.960 2902.510 3490.240 ;
        RECT 2904.530 3489.960 2904.810 3490.240 ;
        RECT 2904.530 3255.360 2904.810 3255.640 ;
        RECT 2904.530 3020.760 2904.810 3021.040 ;
        RECT 2904.530 2786.160 2904.810 2786.440 ;
        RECT 2904.530 2551.560 2904.810 2551.840 ;
        RECT 2904.530 2316.960 2904.810 2317.240 ;
        RECT 2901.310 2082.360 2901.590 2082.640 ;
        RECT 2904.530 2082.360 2904.810 2082.640 ;
        RECT 1986.830 1046.040 1987.110 1046.320 ;
      LAYER met3 ;
        RECT 2902.205 3490.250 2902.535 3490.265 ;
        RECT 2904.505 3490.250 2904.835 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2902.205 3489.950 2924.800 3490.250 ;
        RECT 2902.205 3489.935 2902.535 3489.950 ;
        RECT 2904.505 3489.935 2904.835 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
        RECT 2904.505 3255.650 2904.835 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2904.505 3255.350 2924.800 3255.650 ;
        RECT 2904.505 3255.335 2904.835 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
        RECT 2904.505 3021.050 2904.835 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2904.505 3020.750 2924.800 3021.050 ;
        RECT 2904.505 3020.735 2904.835 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
        RECT 2904.505 2786.450 2904.835 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2904.505 2786.150 2924.800 2786.450 ;
        RECT 2904.505 2786.135 2904.835 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
        RECT 2904.505 2551.850 2904.835 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2904.505 2551.550 2924.800 2551.850 ;
        RECT 2904.505 2551.535 2904.835 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
        RECT 2904.505 2317.250 2904.835 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2904.505 2316.950 2924.800 2317.250 ;
        RECT 2904.505 2316.935 2904.835 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
        RECT 2901.285 2082.650 2901.615 2082.665 ;
        RECT 2904.505 2082.650 2904.835 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2901.285 2082.350 2924.800 2082.650 ;
        RECT 2901.285 2082.335 2901.615 2082.350 ;
        RECT 2904.505 2082.335 2904.835 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
        RECT 1966.720 1046.330 1970.720 1046.520 ;
        RECT 1986.805 1046.330 1987.135 1046.345 ;
        RECT 1966.720 1046.030 1987.135 1046.330 ;
        RECT 1966.720 1045.920 1970.720 1046.030 ;
        RECT 1986.805 1046.015 1987.135 1046.030 ;
    END
  END io_oeb[10]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1897.670 1118.330 1897.950 1120.000 ;
        RECT 1899.430 1118.330 1899.710 1118.445 ;
        RECT 1897.670 1118.190 1899.710 1118.330 ;
        RECT 1897.670 1116.000 1897.950 1118.190 ;
        RECT 1899.430 1118.075 1899.710 1118.190 ;
        RECT 2916.950 16.475 2917.230 16.845 ;
        RECT 2917.020 2.400 2917.160 16.475 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
      LAYER via2 ;
        RECT 1899.430 1118.120 1899.710 1118.400 ;
        RECT 2916.950 16.520 2917.230 16.800 ;
      LAYER met3 ;
        RECT 1899.405 1118.410 1899.735 1118.425 ;
        RECT 1903.750 1118.410 1904.130 1118.420 ;
        RECT 1899.405 1118.110 1904.130 1118.410 ;
        RECT 1899.405 1118.095 1899.735 1118.110 ;
        RECT 1903.750 1118.100 1904.130 1118.110 ;
        RECT 1903.750 16.810 1904.130 16.820 ;
        RECT 2916.925 16.810 2917.255 16.825 ;
        RECT 1903.750 16.510 2917.255 16.810 ;
        RECT 1903.750 16.500 1904.130 16.510 ;
        RECT 2916.925 16.495 2917.255 16.510 ;
      LAYER via3 ;
        RECT 1903.780 1118.100 1904.100 1118.420 ;
        RECT 1903.780 16.500 1904.100 16.820 ;
      LAYER met4 ;
        RECT 1903.775 1118.095 1904.105 1118.425 ;
        RECT 1903.790 16.825 1904.090 1118.095 ;
        RECT 1903.775 16.495 1904.105 16.825 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 40.550 3504.960 40.870 3505.020 ;
        RECT 364.850 3504.960 365.170 3505.020 ;
        RECT 689.150 3504.960 689.470 3505.020 ;
        RECT 1013.910 3504.960 1014.230 3505.020 ;
        RECT 40.550 3504.820 1014.230 3504.960 ;
        RECT 40.550 3504.760 40.870 3504.820 ;
        RECT 364.850 3504.760 365.170 3504.820 ;
        RECT 689.150 3504.760 689.470 3504.820 ;
        RECT 1013.910 3504.760 1014.230 3504.820 ;
        RECT 37.790 3498.500 38.110 3498.560 ;
        RECT 40.550 3498.500 40.870 3498.560 ;
        RECT 37.790 3498.360 40.870 3498.500 ;
        RECT 37.790 3498.300 38.110 3498.360 ;
        RECT 40.550 3498.300 40.870 3498.360 ;
        RECT 16.170 3267.980 16.490 3268.040 ;
        RECT 37.790 3267.980 38.110 3268.040 ;
        RECT 16.170 3267.840 38.110 3267.980 ;
        RECT 16.170 3267.780 16.490 3267.840 ;
        RECT 37.790 3267.780 38.110 3267.840 ;
        RECT 13.870 2121.840 14.190 2121.900 ;
        RECT 16.170 2121.840 16.490 2121.900 ;
        RECT 1472.990 2121.840 1473.310 2121.900 ;
        RECT 13.870 2121.700 1473.310 2121.840 ;
        RECT 13.870 2121.640 14.190 2121.700 ;
        RECT 16.170 2121.640 16.490 2121.700 ;
        RECT 1472.990 2121.640 1473.310 2121.700 ;
        RECT 1472.990 910.420 1473.310 910.480 ;
        RECT 1932.530 910.420 1932.850 910.480 ;
        RECT 1472.990 910.280 1932.850 910.420 ;
        RECT 1472.990 910.220 1473.310 910.280 ;
        RECT 1932.530 910.220 1932.850 910.280 ;
      LAYER via ;
        RECT 40.580 3504.760 40.840 3505.020 ;
        RECT 364.880 3504.760 365.140 3505.020 ;
        RECT 689.180 3504.760 689.440 3505.020 ;
        RECT 1013.940 3504.760 1014.200 3505.020 ;
        RECT 37.820 3498.300 38.080 3498.560 ;
        RECT 40.580 3498.300 40.840 3498.560 ;
        RECT 16.200 3267.780 16.460 3268.040 ;
        RECT 37.820 3267.780 38.080 3268.040 ;
        RECT 13.900 2121.640 14.160 2121.900 ;
        RECT 16.200 2121.640 16.460 2121.900 ;
        RECT 1473.020 2121.640 1473.280 2121.900 ;
        RECT 1473.020 910.220 1473.280 910.480 ;
        RECT 1932.560 910.220 1932.820 910.480 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 40.640 3505.050 40.780 3517.600 ;
        RECT 364.940 3505.050 365.080 3517.600 ;
        RECT 689.240 3505.050 689.380 3517.600 ;
        RECT 1014.000 3505.050 1014.140 3517.600 ;
        RECT 40.580 3504.730 40.840 3505.050 ;
        RECT 364.880 3504.730 365.140 3505.050 ;
        RECT 689.180 3504.730 689.440 3505.050 ;
        RECT 1013.940 3504.730 1014.200 3505.050 ;
        RECT 40.640 3498.590 40.780 3504.730 ;
        RECT 37.820 3498.270 38.080 3498.590 ;
        RECT 40.580 3498.270 40.840 3498.590 ;
        RECT 37.880 3268.070 38.020 3498.270 ;
        RECT 16.200 3267.925 16.460 3268.070 ;
        RECT 13.890 3267.555 14.170 3267.925 ;
        RECT 16.190 3267.555 16.470 3267.925 ;
        RECT 37.820 3267.750 38.080 3268.070 ;
        RECT 13.960 2980.285 14.100 3267.555 ;
        RECT 13.890 2979.915 14.170 2980.285 ;
        RECT 13.960 2693.325 14.100 2979.915 ;
        RECT 13.890 2692.955 14.170 2693.325 ;
        RECT 13.960 2405.685 14.100 2692.955 ;
        RECT 13.890 2405.315 14.170 2405.685 ;
        RECT 13.960 2121.930 14.100 2405.315 ;
        RECT 13.900 2121.610 14.160 2121.930 ;
        RECT 16.200 2121.610 16.460 2121.930 ;
        RECT 1473.020 2121.610 1473.280 2121.930 ;
        RECT 16.260 2118.725 16.400 2121.610 ;
        RECT 16.190 2118.355 16.470 2118.725 ;
        RECT 1473.080 910.510 1473.220 2121.610 ;
        RECT 1932.630 920.380 1932.910 924.000 ;
        RECT 1932.620 920.000 1932.910 920.380 ;
        RECT 1932.620 910.510 1932.760 920.000 ;
        RECT 1473.020 910.190 1473.280 910.510 ;
        RECT 1932.560 910.190 1932.820 910.510 ;
      LAYER via2 ;
        RECT 13.890 3267.600 14.170 3267.880 ;
        RECT 16.190 3267.600 16.470 3267.880 ;
        RECT 13.890 2979.960 14.170 2980.240 ;
        RECT 13.890 2693.000 14.170 2693.280 ;
        RECT 13.890 2405.360 14.170 2405.640 ;
        RECT 16.190 2118.400 16.470 2118.680 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 13.865 3267.890 14.195 3267.905 ;
        RECT 16.165 3267.890 16.495 3267.905 ;
        RECT -4.800 3267.590 16.495 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 13.865 3267.575 14.195 3267.590 ;
        RECT 16.165 3267.575 16.495 3267.590 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 13.865 2980.250 14.195 2980.265 ;
        RECT -4.800 2979.950 14.195 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 13.865 2979.935 14.195 2979.950 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 13.865 2693.290 14.195 2693.305 ;
        RECT -4.800 2692.990 14.195 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 13.865 2692.975 14.195 2692.990 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 13.865 2405.650 14.195 2405.665 ;
        RECT -4.800 2405.350 14.195 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 13.865 2405.335 14.195 2405.350 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 16.165 2118.690 16.495 2118.705 ;
        RECT -4.800 2118.390 16.495 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 16.165 2118.375 16.495 2118.390 ;
    END
  END io_oeb[20]
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.320 7.020 3529.000 ;
        RECT 184.020 -9.320 187.020 3529.000 ;
        RECT 364.020 -9.320 367.020 3529.000 ;
        RECT 544.020 -9.320 547.020 3529.000 ;
        RECT 724.020 -9.320 727.020 3529.000 ;
        RECT 904.020 -9.320 907.020 3529.000 ;
        RECT 1084.020 -9.320 1087.020 3529.000 ;
        RECT 1264.020 -9.320 1267.020 3529.000 ;
        RECT 1444.020 -9.320 1447.020 3529.000 ;
        RECT 1624.020 -9.320 1627.020 3529.000 ;
        RECT 1804.020 -9.320 1807.020 3529.000 ;
        RECT 1984.020 -9.320 1987.020 3529.000 ;
        RECT 2164.020 -9.320 2167.020 3529.000 ;
        RECT 2344.020 -9.320 2347.020 3529.000 ;
        RECT 2524.020 -9.320 2527.020 3529.000 ;
        RECT 2704.020 -9.320 2707.020 3529.000 ;
        RECT 2884.020 -9.320 2887.020 3529.000 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 544.930 2711.090 546.110 2712.270 ;
        RECT 544.930 2709.490 546.110 2710.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 544.930 1991.090 546.110 1992.270 ;
        RECT 544.930 1989.490 546.110 1990.670 ;
        RECT 544.930 1811.090 546.110 1812.270 ;
        RECT 544.930 1809.490 546.110 1810.670 ;
        RECT 544.930 1631.090 546.110 1632.270 ;
        RECT 544.930 1629.490 546.110 1630.670 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 724.930 2171.090 726.110 2172.270 ;
        RECT 724.930 2169.490 726.110 2170.670 ;
        RECT 724.930 1991.090 726.110 1992.270 ;
        RECT 724.930 1989.490 726.110 1990.670 ;
        RECT 724.930 1811.090 726.110 1812.270 ;
        RECT 724.930 1809.490 726.110 1810.670 ;
        RECT 724.930 1631.090 726.110 1632.270 ;
        RECT 724.930 1629.490 726.110 1630.670 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 904.930 2531.090 906.110 2532.270 ;
        RECT 904.930 2529.490 906.110 2530.670 ;
        RECT 904.930 2351.090 906.110 2352.270 ;
        RECT 904.930 2349.490 906.110 2350.670 ;
        RECT 904.930 2171.090 906.110 2172.270 ;
        RECT 904.930 2169.490 906.110 2170.670 ;
        RECT 904.930 1991.090 906.110 1992.270 ;
        RECT 904.930 1989.490 906.110 1990.670 ;
        RECT 904.930 1811.090 906.110 1812.270 ;
        RECT 904.930 1809.490 906.110 1810.670 ;
        RECT 904.930 1631.090 906.110 1632.270 ;
        RECT 904.930 1629.490 906.110 1630.670 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1084.930 2711.090 1086.110 2712.270 ;
        RECT 1084.930 2709.490 1086.110 2710.670 ;
        RECT 1084.930 2531.090 1086.110 2532.270 ;
        RECT 1084.930 2529.490 1086.110 2530.670 ;
        RECT 1084.930 2351.090 1086.110 2352.270 ;
        RECT 1084.930 2349.490 1086.110 2350.670 ;
        RECT 1084.930 2171.090 1086.110 2172.270 ;
        RECT 1084.930 2169.490 1086.110 2170.670 ;
        RECT 1084.930 1991.090 1086.110 1992.270 ;
        RECT 1084.930 1989.490 1086.110 1990.670 ;
        RECT 1084.930 1811.090 1086.110 1812.270 ;
        RECT 1084.930 1809.490 1086.110 1810.670 ;
        RECT 1084.930 1631.090 1086.110 1632.270 ;
        RECT 1084.930 1629.490 1086.110 1630.670 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 1264.930 2711.090 1266.110 2712.270 ;
        RECT 1264.930 2709.490 1266.110 2710.670 ;
        RECT 1264.930 2531.090 1266.110 2532.270 ;
        RECT 1264.930 2529.490 1266.110 2530.670 ;
        RECT 1264.930 2351.090 1266.110 2352.270 ;
        RECT 1264.930 2349.490 1266.110 2350.670 ;
        RECT 1264.930 2171.090 1266.110 2172.270 ;
        RECT 1264.930 2169.490 1266.110 2170.670 ;
        RECT 1264.930 1991.090 1266.110 1992.270 ;
        RECT 1264.930 1989.490 1266.110 1990.670 ;
        RECT 1264.930 1811.090 1266.110 1812.270 ;
        RECT 1264.930 1809.490 1266.110 1810.670 ;
        RECT 1264.930 1631.090 1266.110 1632.270 ;
        RECT 1264.930 1629.490 1266.110 1630.670 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1624.930 2891.090 1626.110 2892.270 ;
        RECT 1624.930 2889.490 1626.110 2890.670 ;
        RECT 1624.930 2711.090 1626.110 2712.270 ;
        RECT 1624.930 2709.490 1626.110 2710.670 ;
        RECT 1624.930 2531.090 1626.110 2532.270 ;
        RECT 1624.930 2529.490 1626.110 2530.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1624.930 1991.090 1626.110 1992.270 ;
        RECT 1624.930 1989.490 1626.110 1990.670 ;
        RECT 1624.930 1811.090 1626.110 1812.270 ;
        RECT 1624.930 1809.490 1626.110 1810.670 ;
        RECT 1624.930 1631.090 1626.110 1632.270 ;
        RECT 1624.930 1629.490 1626.110 1630.670 ;
        RECT 1624.930 1451.090 1626.110 1452.270 ;
        RECT 1624.930 1449.490 1626.110 1450.670 ;
        RECT 1624.930 1271.090 1626.110 1272.270 ;
        RECT 1624.930 1269.490 1626.110 1270.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1624.930 911.090 1626.110 912.270 ;
        RECT 1624.930 909.490 1626.110 910.670 ;
        RECT 1624.930 731.090 1626.110 732.270 ;
        RECT 1624.930 729.490 1626.110 730.670 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1804.930 2891.090 1806.110 2892.270 ;
        RECT 1804.930 2889.490 1806.110 2890.670 ;
        RECT 1804.930 2711.090 1806.110 2712.270 ;
        RECT 1804.930 2709.490 1806.110 2710.670 ;
        RECT 1804.930 2531.090 1806.110 2532.270 ;
        RECT 1804.930 2529.490 1806.110 2530.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1804.930 1991.090 1806.110 1992.270 ;
        RECT 1804.930 1989.490 1806.110 1990.670 ;
        RECT 1804.930 1811.090 1806.110 1812.270 ;
        RECT 1804.930 1809.490 1806.110 1810.670 ;
        RECT 1804.930 1631.090 1806.110 1632.270 ;
        RECT 1804.930 1629.490 1806.110 1630.670 ;
        RECT 1804.930 1451.090 1806.110 1452.270 ;
        RECT 1804.930 1449.490 1806.110 1450.670 ;
        RECT 1804.930 1271.090 1806.110 1272.270 ;
        RECT 1804.930 1269.490 1806.110 1270.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1804.930 911.090 1806.110 912.270 ;
        RECT 1804.930 909.490 1806.110 910.670 ;
        RECT 1804.930 731.090 1806.110 732.270 ;
        RECT 1804.930 729.490 1806.110 730.670 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 1984.930 1991.090 1986.110 1992.270 ;
        RECT 1984.930 1989.490 1986.110 1990.670 ;
        RECT 1984.930 1811.090 1986.110 1812.270 ;
        RECT 1984.930 1809.490 1986.110 1810.670 ;
        RECT 1984.930 1631.090 1986.110 1632.270 ;
        RECT 1984.930 1629.490 1986.110 1630.670 ;
        RECT 1984.930 1451.090 1986.110 1452.270 ;
        RECT 1984.930 1449.490 1986.110 1450.670 ;
        RECT 1984.930 1271.090 1986.110 1272.270 ;
        RECT 1984.930 1269.490 1986.110 1270.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 1984.930 911.090 1986.110 912.270 ;
        RECT 1984.930 909.490 1986.110 910.670 ;
        RECT 1984.930 731.090 1986.110 732.270 ;
        RECT 1984.930 729.490 1986.110 730.670 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2164.930 1451.090 2166.110 1452.270 ;
        RECT 2164.930 1449.490 2166.110 1450.670 ;
        RECT 2164.930 1271.090 2166.110 1272.270 ;
        RECT 2164.930 1269.490 2166.110 1270.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2164.930 911.090 2166.110 912.270 ;
        RECT 2164.930 909.490 2166.110 910.670 ;
        RECT 2164.930 731.090 2166.110 732.270 ;
        RECT 2164.930 729.490 2166.110 730.670 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2344.930 1811.090 2346.110 1812.270 ;
        RECT 2344.930 1809.490 2346.110 1810.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.680 3429.380 2934.300 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.680 3249.380 2934.300 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.680 3069.380 2934.300 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 544.020 2892.380 547.020 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1084.020 2892.380 1087.020 2892.390 ;
        RECT 1264.020 2892.380 1267.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1624.020 2892.380 1627.020 2892.390 ;
        RECT 1804.020 2892.380 1807.020 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2344.020 2892.380 2347.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.680 2889.380 2934.300 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 544.020 2889.370 547.020 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1084.020 2889.370 1087.020 2889.380 ;
        RECT 1264.020 2889.370 1267.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1624.020 2889.370 1627.020 2889.380 ;
        RECT 1804.020 2889.370 1807.020 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2344.020 2889.370 2347.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 544.020 2712.380 547.020 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 904.020 2712.380 907.020 2712.390 ;
        RECT 1084.020 2712.380 1087.020 2712.390 ;
        RECT 1264.020 2712.380 1267.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1624.020 2712.380 1627.020 2712.390 ;
        RECT 1804.020 2712.380 1807.020 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.680 2709.380 2934.300 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 544.020 2709.370 547.020 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 904.020 2709.370 907.020 2709.380 ;
        RECT 1084.020 2709.370 1087.020 2709.380 ;
        RECT 1264.020 2709.370 1267.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1624.020 2709.370 1627.020 2709.380 ;
        RECT 1804.020 2709.370 1807.020 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 544.020 2532.380 547.020 2532.390 ;
        RECT 724.020 2532.380 727.020 2532.390 ;
        RECT 904.020 2532.380 907.020 2532.390 ;
        RECT 1084.020 2532.380 1087.020 2532.390 ;
        RECT 1264.020 2532.380 1267.020 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1624.020 2532.380 1627.020 2532.390 ;
        RECT 1804.020 2532.380 1807.020 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.680 2529.380 2934.300 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 544.020 2529.370 547.020 2529.380 ;
        RECT 724.020 2529.370 727.020 2529.380 ;
        RECT 904.020 2529.370 907.020 2529.380 ;
        RECT 1084.020 2529.370 1087.020 2529.380 ;
        RECT 1264.020 2529.370 1267.020 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1624.020 2529.370 1627.020 2529.380 ;
        RECT 1804.020 2529.370 1807.020 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 544.020 2352.380 547.020 2352.390 ;
        RECT 724.020 2352.380 727.020 2352.390 ;
        RECT 904.020 2352.380 907.020 2352.390 ;
        RECT 1084.020 2352.380 1087.020 2352.390 ;
        RECT 1264.020 2352.380 1267.020 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1624.020 2352.380 1627.020 2352.390 ;
        RECT 1804.020 2352.380 1807.020 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.680 2349.380 2934.300 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 544.020 2349.370 547.020 2349.380 ;
        RECT 724.020 2349.370 727.020 2349.380 ;
        RECT 904.020 2349.370 907.020 2349.380 ;
        RECT 1084.020 2349.370 1087.020 2349.380 ;
        RECT 1264.020 2349.370 1267.020 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1624.020 2349.370 1627.020 2349.380 ;
        RECT 1804.020 2349.370 1807.020 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 544.020 2172.380 547.020 2172.390 ;
        RECT 724.020 2172.380 727.020 2172.390 ;
        RECT 904.020 2172.380 907.020 2172.390 ;
        RECT 1084.020 2172.380 1087.020 2172.390 ;
        RECT 1264.020 2172.380 1267.020 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.680 2169.380 2934.300 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 544.020 2169.370 547.020 2169.380 ;
        RECT 724.020 2169.370 727.020 2169.380 ;
        RECT 904.020 2169.370 907.020 2169.380 ;
        RECT 1084.020 2169.370 1087.020 2169.380 ;
        RECT 1264.020 2169.370 1267.020 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 544.020 1992.380 547.020 1992.390 ;
        RECT 724.020 1992.380 727.020 1992.390 ;
        RECT 904.020 1992.380 907.020 1992.390 ;
        RECT 1084.020 1992.380 1087.020 1992.390 ;
        RECT 1264.020 1992.380 1267.020 1992.390 ;
        RECT 1444.020 1992.380 1447.020 1992.390 ;
        RECT 1624.020 1992.380 1627.020 1992.390 ;
        RECT 1804.020 1992.380 1807.020 1992.390 ;
        RECT 1984.020 1992.380 1987.020 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.680 1989.380 2934.300 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 544.020 1989.370 547.020 1989.380 ;
        RECT 724.020 1989.370 727.020 1989.380 ;
        RECT 904.020 1989.370 907.020 1989.380 ;
        RECT 1084.020 1989.370 1087.020 1989.380 ;
        RECT 1264.020 1989.370 1267.020 1989.380 ;
        RECT 1444.020 1989.370 1447.020 1989.380 ;
        RECT 1624.020 1989.370 1627.020 1989.380 ;
        RECT 1804.020 1989.370 1807.020 1989.380 ;
        RECT 1984.020 1989.370 1987.020 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 364.020 1812.380 367.020 1812.390 ;
        RECT 544.020 1812.380 547.020 1812.390 ;
        RECT 724.020 1812.380 727.020 1812.390 ;
        RECT 904.020 1812.380 907.020 1812.390 ;
        RECT 1084.020 1812.380 1087.020 1812.390 ;
        RECT 1264.020 1812.380 1267.020 1812.390 ;
        RECT 1444.020 1812.380 1447.020 1812.390 ;
        RECT 1624.020 1812.380 1627.020 1812.390 ;
        RECT 1804.020 1812.380 1807.020 1812.390 ;
        RECT 1984.020 1812.380 1987.020 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2344.020 1812.380 2347.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.680 1809.380 2934.300 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 364.020 1809.370 367.020 1809.380 ;
        RECT 544.020 1809.370 547.020 1809.380 ;
        RECT 724.020 1809.370 727.020 1809.380 ;
        RECT 904.020 1809.370 907.020 1809.380 ;
        RECT 1084.020 1809.370 1087.020 1809.380 ;
        RECT 1264.020 1809.370 1267.020 1809.380 ;
        RECT 1444.020 1809.370 1447.020 1809.380 ;
        RECT 1624.020 1809.370 1627.020 1809.380 ;
        RECT 1804.020 1809.370 1807.020 1809.380 ;
        RECT 1984.020 1809.370 1987.020 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2344.020 1809.370 2347.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 544.020 1632.380 547.020 1632.390 ;
        RECT 724.020 1632.380 727.020 1632.390 ;
        RECT 904.020 1632.380 907.020 1632.390 ;
        RECT 1084.020 1632.380 1087.020 1632.390 ;
        RECT 1264.020 1632.380 1267.020 1632.390 ;
        RECT 1444.020 1632.380 1447.020 1632.390 ;
        RECT 1624.020 1632.380 1627.020 1632.390 ;
        RECT 1804.020 1632.380 1807.020 1632.390 ;
        RECT 1984.020 1632.380 1987.020 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.680 1629.380 2934.300 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 544.020 1629.370 547.020 1629.380 ;
        RECT 724.020 1629.370 727.020 1629.380 ;
        RECT 904.020 1629.370 907.020 1629.380 ;
        RECT 1084.020 1629.370 1087.020 1629.380 ;
        RECT 1264.020 1629.370 1267.020 1629.380 ;
        RECT 1444.020 1629.370 1447.020 1629.380 ;
        RECT 1624.020 1629.370 1627.020 1629.380 ;
        RECT 1804.020 1629.370 1807.020 1629.380 ;
        RECT 1984.020 1629.370 1987.020 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1444.020 1452.380 1447.020 1452.390 ;
        RECT 1624.020 1452.380 1627.020 1452.390 ;
        RECT 1804.020 1452.380 1807.020 1452.390 ;
        RECT 1984.020 1452.380 1987.020 1452.390 ;
        RECT 2164.020 1452.380 2167.020 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.680 1449.380 2934.300 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1444.020 1449.370 1447.020 1449.380 ;
        RECT 1624.020 1449.370 1627.020 1449.380 ;
        RECT 1804.020 1449.370 1807.020 1449.380 ;
        RECT 1984.020 1449.370 1987.020 1449.380 ;
        RECT 2164.020 1449.370 2167.020 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1444.020 1272.380 1447.020 1272.390 ;
        RECT 1624.020 1272.380 1627.020 1272.390 ;
        RECT 1804.020 1272.380 1807.020 1272.390 ;
        RECT 1984.020 1272.380 1987.020 1272.390 ;
        RECT 2164.020 1272.380 2167.020 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.680 1269.380 2934.300 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1444.020 1269.370 1447.020 1269.380 ;
        RECT 1624.020 1269.370 1627.020 1269.380 ;
        RECT 1804.020 1269.370 1807.020 1269.380 ;
        RECT 1984.020 1269.370 1987.020 1269.380 ;
        RECT 2164.020 1269.370 2167.020 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.680 1089.380 2934.300 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1624.020 912.380 1627.020 912.390 ;
        RECT 1804.020 912.380 1807.020 912.390 ;
        RECT 1984.020 912.380 1987.020 912.390 ;
        RECT 2164.020 912.380 2167.020 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.680 909.380 2934.300 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1624.020 909.370 1627.020 909.380 ;
        RECT 1804.020 909.370 1807.020 909.380 ;
        RECT 1984.020 909.370 1987.020 909.380 ;
        RECT 2164.020 909.370 2167.020 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1624.020 732.380 1627.020 732.390 ;
        RECT 1804.020 732.380 1807.020 732.390 ;
        RECT 1984.020 732.380 1987.020 732.390 ;
        RECT 2164.020 732.380 2167.020 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.680 729.380 2934.300 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1624.020 729.370 1627.020 729.380 ;
        RECT 1804.020 729.370 1807.020 729.380 ;
        RECT 1984.020 729.370 1987.020 729.380 ;
        RECT 2164.020 729.370 2167.020 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1624.020 552.380 1627.020 552.390 ;
        RECT 1804.020 552.380 1807.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.680 549.380 2934.300 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1624.020 549.370 1627.020 549.380 ;
        RECT 1804.020 549.370 1807.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.680 369.380 2934.300 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.680 189.380 2934.300 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.680 9.380 2934.300 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 -9.320 97.020 3529.000 ;
        RECT 274.020 -9.320 277.020 3529.000 ;
        RECT 454.020 -9.320 457.020 3529.000 ;
        RECT 634.020 -9.320 637.020 3529.000 ;
        RECT 814.020 -9.320 817.020 3529.000 ;
        RECT 994.020 -9.320 997.020 3529.000 ;
        RECT 1174.020 -9.320 1177.020 3529.000 ;
        RECT 1354.020 -9.320 1357.020 3529.000 ;
        RECT 1534.020 -9.320 1537.020 3529.000 ;
        RECT 1714.020 -9.320 1717.020 3529.000 ;
        RECT 1894.020 -9.320 1897.020 3529.000 ;
        RECT 2074.020 -9.320 2077.020 3529.000 ;
        RECT 2254.020 -9.320 2257.020 3529.000 ;
        RECT 2434.020 -9.320 2437.020 3529.000 ;
        RECT 2614.020 -9.320 2617.020 3529.000 ;
        RECT 2794.020 -9.320 2797.020 3529.000 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER via4 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT -13.770 3341.090 -12.590 3342.270 ;
        RECT -13.770 3339.490 -12.590 3340.670 ;
        RECT -13.770 3161.090 -12.590 3162.270 ;
        RECT -13.770 3159.490 -12.590 3160.670 ;
        RECT -13.770 2981.090 -12.590 2982.270 ;
        RECT -13.770 2979.490 -12.590 2980.670 ;
        RECT -13.770 2801.090 -12.590 2802.270 ;
        RECT -13.770 2799.490 -12.590 2800.670 ;
        RECT -13.770 2621.090 -12.590 2622.270 ;
        RECT -13.770 2619.490 -12.590 2620.670 ;
        RECT -13.770 2441.090 -12.590 2442.270 ;
        RECT -13.770 2439.490 -12.590 2440.670 ;
        RECT -13.770 2261.090 -12.590 2262.270 ;
        RECT -13.770 2259.490 -12.590 2260.670 ;
        RECT -13.770 2081.090 -12.590 2082.270 ;
        RECT -13.770 2079.490 -12.590 2080.670 ;
        RECT -13.770 1901.090 -12.590 1902.270 ;
        RECT -13.770 1899.490 -12.590 1900.670 ;
        RECT -13.770 1721.090 -12.590 1722.270 ;
        RECT -13.770 1719.490 -12.590 1720.670 ;
        RECT -13.770 1541.090 -12.590 1542.270 ;
        RECT -13.770 1539.490 -12.590 1540.670 ;
        RECT -13.770 1361.090 -12.590 1362.270 ;
        RECT -13.770 1359.490 -12.590 1360.670 ;
        RECT -13.770 1181.090 -12.590 1182.270 ;
        RECT -13.770 1179.490 -12.590 1180.670 ;
        RECT -13.770 1001.090 -12.590 1002.270 ;
        RECT -13.770 999.490 -12.590 1000.670 ;
        RECT -13.770 821.090 -12.590 822.270 ;
        RECT -13.770 819.490 -12.590 820.670 ;
        RECT -13.770 641.090 -12.590 642.270 ;
        RECT -13.770 639.490 -12.590 640.670 ;
        RECT -13.770 461.090 -12.590 462.270 ;
        RECT -13.770 459.490 -12.590 460.670 ;
        RECT -13.770 281.090 -12.590 282.270 ;
        RECT -13.770 279.490 -12.590 280.670 ;
        RECT -13.770 101.090 -12.590 102.270 ;
        RECT -13.770 99.490 -12.590 100.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 454.930 2621.090 456.110 2622.270 ;
        RECT 454.930 2619.490 456.110 2620.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 454.930 2081.090 456.110 2082.270 ;
        RECT 454.930 2079.490 456.110 2080.670 ;
        RECT 454.930 1901.090 456.110 1902.270 ;
        RECT 454.930 1899.490 456.110 1900.670 ;
        RECT 454.930 1721.090 456.110 1722.270 ;
        RECT 454.930 1719.490 456.110 1720.670 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 634.930 2081.090 636.110 2082.270 ;
        RECT 634.930 2079.490 636.110 2080.670 ;
        RECT 634.930 1901.090 636.110 1902.270 ;
        RECT 634.930 1899.490 636.110 1900.670 ;
        RECT 634.930 1721.090 636.110 1722.270 ;
        RECT 634.930 1719.490 636.110 1720.670 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 814.930 2441.090 816.110 2442.270 ;
        RECT 814.930 2439.490 816.110 2440.670 ;
        RECT 814.930 2261.090 816.110 2262.270 ;
        RECT 814.930 2259.490 816.110 2260.670 ;
        RECT 814.930 2081.090 816.110 2082.270 ;
        RECT 814.930 2079.490 816.110 2080.670 ;
        RECT 814.930 1901.090 816.110 1902.270 ;
        RECT 814.930 1899.490 816.110 1900.670 ;
        RECT 814.930 1721.090 816.110 1722.270 ;
        RECT 814.930 1719.490 816.110 1720.670 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 814.930 1001.090 816.110 1002.270 ;
        RECT 814.930 999.490 816.110 1000.670 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 994.930 2621.090 996.110 2622.270 ;
        RECT 994.930 2619.490 996.110 2620.670 ;
        RECT 994.930 2441.090 996.110 2442.270 ;
        RECT 994.930 2439.490 996.110 2440.670 ;
        RECT 994.930 2261.090 996.110 2262.270 ;
        RECT 994.930 2259.490 996.110 2260.670 ;
        RECT 994.930 2081.090 996.110 2082.270 ;
        RECT 994.930 2079.490 996.110 2080.670 ;
        RECT 994.930 1901.090 996.110 1902.270 ;
        RECT 994.930 1899.490 996.110 1900.670 ;
        RECT 994.930 1721.090 996.110 1722.270 ;
        RECT 994.930 1719.490 996.110 1720.670 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 994.930 1001.090 996.110 1002.270 ;
        RECT 994.930 999.490 996.110 1000.670 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 1174.930 2621.090 1176.110 2622.270 ;
        RECT 1174.930 2619.490 1176.110 2620.670 ;
        RECT 1174.930 2441.090 1176.110 2442.270 ;
        RECT 1174.930 2439.490 1176.110 2440.670 ;
        RECT 1174.930 2261.090 1176.110 2262.270 ;
        RECT 1174.930 2259.490 1176.110 2260.670 ;
        RECT 1174.930 2081.090 1176.110 2082.270 ;
        RECT 1174.930 2079.490 1176.110 2080.670 ;
        RECT 1174.930 1901.090 1176.110 1902.270 ;
        RECT 1174.930 1899.490 1176.110 1900.670 ;
        RECT 1174.930 1721.090 1176.110 1722.270 ;
        RECT 1174.930 1719.490 1176.110 1720.670 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1174.930 1001.090 1176.110 1002.270 ;
        RECT 1174.930 999.490 1176.110 1000.670 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1354.930 2441.090 1356.110 2442.270 ;
        RECT 1354.930 2439.490 1356.110 2440.670 ;
        RECT 1354.930 2261.090 1356.110 2262.270 ;
        RECT 1354.930 2259.490 1356.110 2260.670 ;
        RECT 1354.930 2081.090 1356.110 2082.270 ;
        RECT 1354.930 2079.490 1356.110 2080.670 ;
        RECT 1354.930 1901.090 1356.110 1902.270 ;
        RECT 1354.930 1899.490 1356.110 1900.670 ;
        RECT 1354.930 1721.090 1356.110 1722.270 ;
        RECT 1354.930 1719.490 1356.110 1720.670 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1354.930 1001.090 1356.110 1002.270 ;
        RECT 1354.930 999.490 1356.110 1000.670 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1534.930 2981.090 1536.110 2982.270 ;
        RECT 1534.930 2979.490 1536.110 2980.670 ;
        RECT 1534.930 2801.090 1536.110 2802.270 ;
        RECT 1534.930 2799.490 1536.110 2800.670 ;
        RECT 1534.930 2621.090 1536.110 2622.270 ;
        RECT 1534.930 2619.490 1536.110 2620.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1534.930 1901.090 1536.110 1902.270 ;
        RECT 1534.930 1899.490 1536.110 1900.670 ;
        RECT 1534.930 1721.090 1536.110 1722.270 ;
        RECT 1534.930 1719.490 1536.110 1720.670 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1534.930 1361.090 1536.110 1362.270 ;
        RECT 1534.930 1359.490 1536.110 1360.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1534.930 1001.090 1536.110 1002.270 ;
        RECT 1534.930 999.490 1536.110 1000.670 ;
        RECT 1534.930 821.090 1536.110 822.270 ;
        RECT 1534.930 819.490 1536.110 820.670 ;
        RECT 1534.930 641.090 1536.110 642.270 ;
        RECT 1534.930 639.490 1536.110 640.670 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1714.930 2981.090 1716.110 2982.270 ;
        RECT 1714.930 2979.490 1716.110 2980.670 ;
        RECT 1714.930 2801.090 1716.110 2802.270 ;
        RECT 1714.930 2799.490 1716.110 2800.670 ;
        RECT 1714.930 2621.090 1716.110 2622.270 ;
        RECT 1714.930 2619.490 1716.110 2620.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1714.930 1901.090 1716.110 1902.270 ;
        RECT 1714.930 1899.490 1716.110 1900.670 ;
        RECT 1714.930 1721.090 1716.110 1722.270 ;
        RECT 1714.930 1719.490 1716.110 1720.670 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1714.930 1361.090 1716.110 1362.270 ;
        RECT 1714.930 1359.490 1716.110 1360.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1714.930 1001.090 1716.110 1002.270 ;
        RECT 1714.930 999.490 1716.110 1000.670 ;
        RECT 1714.930 821.090 1716.110 822.270 ;
        RECT 1714.930 819.490 1716.110 820.670 ;
        RECT 1714.930 641.090 1716.110 642.270 ;
        RECT 1714.930 639.490 1716.110 640.670 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 1894.930 2981.090 1896.110 2982.270 ;
        RECT 1894.930 2979.490 1896.110 2980.670 ;
        RECT 1894.930 2801.090 1896.110 2802.270 ;
        RECT 1894.930 2799.490 1896.110 2800.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 1894.930 1901.090 1896.110 1902.270 ;
        RECT 1894.930 1899.490 1896.110 1900.670 ;
        RECT 1894.930 1721.090 1896.110 1722.270 ;
        RECT 1894.930 1719.490 1896.110 1720.670 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1894.930 1361.090 1896.110 1362.270 ;
        RECT 1894.930 1359.490 1896.110 1360.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 1894.930 1001.090 1896.110 1002.270 ;
        RECT 1894.930 999.490 1896.110 1000.670 ;
        RECT 1894.930 821.090 1896.110 822.270 ;
        RECT 1894.930 819.490 1896.110 820.670 ;
        RECT 1894.930 641.090 1896.110 642.270 ;
        RECT 1894.930 639.490 1896.110 640.670 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 2074.930 1901.090 2076.110 1902.270 ;
        RECT 2074.930 1899.490 2076.110 1900.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2074.930 1361.090 2076.110 1362.270 ;
        RECT 2074.930 1359.490 2076.110 1360.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2074.930 1001.090 2076.110 1002.270 ;
        RECT 2074.930 999.490 2076.110 1000.670 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2434.930 1901.090 2436.110 1902.270 ;
        RECT 2434.930 1899.490 2436.110 1900.670 ;
        RECT 2434.930 1721.090 2436.110 1722.270 ;
        RECT 2434.930 1719.490 2436.110 1720.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT 2932.210 3341.090 2933.390 3342.270 ;
        RECT 2932.210 3339.490 2933.390 3340.670 ;
        RECT 2932.210 3161.090 2933.390 3162.270 ;
        RECT 2932.210 3159.490 2933.390 3160.670 ;
        RECT 2932.210 2981.090 2933.390 2982.270 ;
        RECT 2932.210 2979.490 2933.390 2980.670 ;
        RECT 2932.210 2801.090 2933.390 2802.270 ;
        RECT 2932.210 2799.490 2933.390 2800.670 ;
        RECT 2932.210 2621.090 2933.390 2622.270 ;
        RECT 2932.210 2619.490 2933.390 2620.670 ;
        RECT 2932.210 2441.090 2933.390 2442.270 ;
        RECT 2932.210 2439.490 2933.390 2440.670 ;
        RECT 2932.210 2261.090 2933.390 2262.270 ;
        RECT 2932.210 2259.490 2933.390 2260.670 ;
        RECT 2932.210 2081.090 2933.390 2082.270 ;
        RECT 2932.210 2079.490 2933.390 2080.670 ;
        RECT 2932.210 1901.090 2933.390 1902.270 ;
        RECT 2932.210 1899.490 2933.390 1900.670 ;
        RECT 2932.210 1721.090 2933.390 1722.270 ;
        RECT 2932.210 1719.490 2933.390 1720.670 ;
        RECT 2932.210 1541.090 2933.390 1542.270 ;
        RECT 2932.210 1539.490 2933.390 1540.670 ;
        RECT 2932.210 1361.090 2933.390 1362.270 ;
        RECT 2932.210 1359.490 2933.390 1360.670 ;
        RECT 2932.210 1181.090 2933.390 1182.270 ;
        RECT 2932.210 1179.490 2933.390 1180.670 ;
        RECT 2932.210 1001.090 2933.390 1002.270 ;
        RECT 2932.210 999.490 2933.390 1000.670 ;
        RECT 2932.210 821.090 2933.390 822.270 ;
        RECT 2932.210 819.490 2933.390 820.670 ;
        RECT 2932.210 641.090 2933.390 642.270 ;
        RECT 2932.210 639.490 2933.390 640.670 ;
        RECT 2932.210 461.090 2933.390 462.270 ;
        RECT 2932.210 459.490 2933.390 460.670 ;
        RECT 2932.210 281.090 2933.390 282.270 ;
        RECT 2932.210 279.490 2933.390 280.670 ;
        RECT 2932.210 101.090 2933.390 102.270 ;
        RECT 2932.210 99.490 2933.390 100.670 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.300 3342.380 2934.300 3342.390 ;
        RECT -14.680 3339.380 2934.300 3342.380 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.300 3339.370 2934.300 3339.380 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.300 3162.380 2934.300 3162.390 ;
        RECT -14.680 3159.380 2934.300 3162.380 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.300 3159.370 2934.300 3159.380 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 454.020 2982.380 457.020 2982.390 ;
        RECT 634.020 2982.380 637.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 994.020 2982.380 997.020 2982.390 ;
        RECT 1174.020 2982.380 1177.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1534.020 2982.380 1537.020 2982.390 ;
        RECT 1714.020 2982.380 1717.020 2982.390 ;
        RECT 1894.020 2982.380 1897.020 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2254.020 2982.380 2257.020 2982.390 ;
        RECT 2434.020 2982.380 2437.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.300 2982.380 2934.300 2982.390 ;
        RECT -14.680 2979.380 2934.300 2982.380 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 454.020 2979.370 457.020 2979.380 ;
        RECT 634.020 2979.370 637.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 994.020 2979.370 997.020 2979.380 ;
        RECT 1174.020 2979.370 1177.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1534.020 2979.370 1537.020 2979.380 ;
        RECT 1714.020 2979.370 1717.020 2979.380 ;
        RECT 1894.020 2979.370 1897.020 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2254.020 2979.370 2257.020 2979.380 ;
        RECT 2434.020 2979.370 2437.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.300 2979.370 2934.300 2979.380 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1534.020 2802.380 1537.020 2802.390 ;
        RECT 1714.020 2802.380 1717.020 2802.390 ;
        RECT 1894.020 2802.380 1897.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2254.020 2802.380 2257.020 2802.390 ;
        RECT 2434.020 2802.380 2437.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.300 2802.380 2934.300 2802.390 ;
        RECT -14.680 2799.380 2934.300 2802.380 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1534.020 2799.370 1537.020 2799.380 ;
        RECT 1714.020 2799.370 1717.020 2799.380 ;
        RECT 1894.020 2799.370 1897.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2254.020 2799.370 2257.020 2799.380 ;
        RECT 2434.020 2799.370 2437.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.300 2799.370 2934.300 2799.380 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 454.020 2622.380 457.020 2622.390 ;
        RECT 634.020 2622.380 637.020 2622.390 ;
        RECT 814.020 2622.380 817.020 2622.390 ;
        RECT 994.020 2622.380 997.020 2622.390 ;
        RECT 1174.020 2622.380 1177.020 2622.390 ;
        RECT 1354.020 2622.380 1357.020 2622.390 ;
        RECT 1534.020 2622.380 1537.020 2622.390 ;
        RECT 1714.020 2622.380 1717.020 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2434.020 2622.380 2437.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.300 2622.380 2934.300 2622.390 ;
        RECT -14.680 2619.380 2934.300 2622.380 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 454.020 2619.370 457.020 2619.380 ;
        RECT 634.020 2619.370 637.020 2619.380 ;
        RECT 814.020 2619.370 817.020 2619.380 ;
        RECT 994.020 2619.370 997.020 2619.380 ;
        RECT 1174.020 2619.370 1177.020 2619.380 ;
        RECT 1354.020 2619.370 1357.020 2619.380 ;
        RECT 1534.020 2619.370 1537.020 2619.380 ;
        RECT 1714.020 2619.370 1717.020 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2434.020 2619.370 2437.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.300 2619.370 2934.300 2619.380 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 454.020 2442.380 457.020 2442.390 ;
        RECT 634.020 2442.380 637.020 2442.390 ;
        RECT 814.020 2442.380 817.020 2442.390 ;
        RECT 994.020 2442.380 997.020 2442.390 ;
        RECT 1174.020 2442.380 1177.020 2442.390 ;
        RECT 1354.020 2442.380 1357.020 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.300 2442.380 2934.300 2442.390 ;
        RECT -14.680 2439.380 2934.300 2442.380 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 454.020 2439.370 457.020 2439.380 ;
        RECT 634.020 2439.370 637.020 2439.380 ;
        RECT 814.020 2439.370 817.020 2439.380 ;
        RECT 994.020 2439.370 997.020 2439.380 ;
        RECT 1174.020 2439.370 1177.020 2439.380 ;
        RECT 1354.020 2439.370 1357.020 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.300 2439.370 2934.300 2439.380 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 814.020 2262.380 817.020 2262.390 ;
        RECT 994.020 2262.380 997.020 2262.390 ;
        RECT 1174.020 2262.380 1177.020 2262.390 ;
        RECT 1354.020 2262.380 1357.020 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.300 2262.380 2934.300 2262.390 ;
        RECT -14.680 2259.380 2934.300 2262.380 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 814.020 2259.370 817.020 2259.380 ;
        RECT 994.020 2259.370 997.020 2259.380 ;
        RECT 1174.020 2259.370 1177.020 2259.380 ;
        RECT 1354.020 2259.370 1357.020 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.300 2259.370 2934.300 2259.380 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 454.020 2082.380 457.020 2082.390 ;
        RECT 634.020 2082.380 637.020 2082.390 ;
        RECT 814.020 2082.380 817.020 2082.390 ;
        RECT 994.020 2082.380 997.020 2082.390 ;
        RECT 1174.020 2082.380 1177.020 2082.390 ;
        RECT 1354.020 2082.380 1357.020 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.300 2082.380 2934.300 2082.390 ;
        RECT -14.680 2079.380 2934.300 2082.380 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 454.020 2079.370 457.020 2079.380 ;
        RECT 634.020 2079.370 637.020 2079.380 ;
        RECT 814.020 2079.370 817.020 2079.380 ;
        RECT 994.020 2079.370 997.020 2079.380 ;
        RECT 1174.020 2079.370 1177.020 2079.380 ;
        RECT 1354.020 2079.370 1357.020 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.300 2079.370 2934.300 2079.380 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 454.020 1902.380 457.020 1902.390 ;
        RECT 634.020 1902.380 637.020 1902.390 ;
        RECT 814.020 1902.380 817.020 1902.390 ;
        RECT 994.020 1902.380 997.020 1902.390 ;
        RECT 1174.020 1902.380 1177.020 1902.390 ;
        RECT 1354.020 1902.380 1357.020 1902.390 ;
        RECT 1534.020 1902.380 1537.020 1902.390 ;
        RECT 1714.020 1902.380 1717.020 1902.390 ;
        RECT 1894.020 1902.380 1897.020 1902.390 ;
        RECT 2074.020 1902.380 2077.020 1902.390 ;
        RECT 2254.020 1902.380 2257.020 1902.390 ;
        RECT 2434.020 1902.380 2437.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.300 1902.380 2934.300 1902.390 ;
        RECT -14.680 1899.380 2934.300 1902.380 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 454.020 1899.370 457.020 1899.380 ;
        RECT 634.020 1899.370 637.020 1899.380 ;
        RECT 814.020 1899.370 817.020 1899.380 ;
        RECT 994.020 1899.370 997.020 1899.380 ;
        RECT 1174.020 1899.370 1177.020 1899.380 ;
        RECT 1354.020 1899.370 1357.020 1899.380 ;
        RECT 1534.020 1899.370 1537.020 1899.380 ;
        RECT 1714.020 1899.370 1717.020 1899.380 ;
        RECT 1894.020 1899.370 1897.020 1899.380 ;
        RECT 2074.020 1899.370 2077.020 1899.380 ;
        RECT 2254.020 1899.370 2257.020 1899.380 ;
        RECT 2434.020 1899.370 2437.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.300 1899.370 2934.300 1899.380 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 454.020 1722.380 457.020 1722.390 ;
        RECT 634.020 1722.380 637.020 1722.390 ;
        RECT 814.020 1722.380 817.020 1722.390 ;
        RECT 994.020 1722.380 997.020 1722.390 ;
        RECT 1174.020 1722.380 1177.020 1722.390 ;
        RECT 1354.020 1722.380 1357.020 1722.390 ;
        RECT 1534.020 1722.380 1537.020 1722.390 ;
        RECT 1714.020 1722.380 1717.020 1722.390 ;
        RECT 1894.020 1722.380 1897.020 1722.390 ;
        RECT 2074.020 1722.380 2077.020 1722.390 ;
        RECT 2254.020 1722.380 2257.020 1722.390 ;
        RECT 2434.020 1722.380 2437.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.300 1722.380 2934.300 1722.390 ;
        RECT -14.680 1719.380 2934.300 1722.380 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 454.020 1719.370 457.020 1719.380 ;
        RECT 634.020 1719.370 637.020 1719.380 ;
        RECT 814.020 1719.370 817.020 1719.380 ;
        RECT 994.020 1719.370 997.020 1719.380 ;
        RECT 1174.020 1719.370 1177.020 1719.380 ;
        RECT 1354.020 1719.370 1357.020 1719.380 ;
        RECT 1534.020 1719.370 1537.020 1719.380 ;
        RECT 1714.020 1719.370 1717.020 1719.380 ;
        RECT 1894.020 1719.370 1897.020 1719.380 ;
        RECT 2074.020 1719.370 2077.020 1719.380 ;
        RECT 2254.020 1719.370 2257.020 1719.380 ;
        RECT 2434.020 1719.370 2437.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.300 1719.370 2934.300 1719.380 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1354.020 1542.380 1357.020 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.300 1542.380 2934.300 1542.390 ;
        RECT -14.680 1539.380 2934.300 1542.380 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1354.020 1539.370 1357.020 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.300 1539.370 2934.300 1539.380 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1534.020 1362.380 1537.020 1362.390 ;
        RECT 1714.020 1362.380 1717.020 1362.390 ;
        RECT 1894.020 1362.380 1897.020 1362.390 ;
        RECT 2074.020 1362.380 2077.020 1362.390 ;
        RECT 2254.020 1362.380 2257.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.300 1362.380 2934.300 1362.390 ;
        RECT -14.680 1359.380 2934.300 1362.380 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1534.020 1359.370 1537.020 1359.380 ;
        RECT 1714.020 1359.370 1717.020 1359.380 ;
        RECT 1894.020 1359.370 1897.020 1359.380 ;
        RECT 2074.020 1359.370 2077.020 1359.380 ;
        RECT 2254.020 1359.370 2257.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.300 1359.370 2934.300 1359.380 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.300 1182.380 2934.300 1182.390 ;
        RECT -14.680 1179.380 2934.300 1182.380 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.300 1179.370 2934.300 1179.380 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 814.020 1002.380 817.020 1002.390 ;
        RECT 994.020 1002.380 997.020 1002.390 ;
        RECT 1174.020 1002.380 1177.020 1002.390 ;
        RECT 1354.020 1002.380 1357.020 1002.390 ;
        RECT 1534.020 1002.380 1537.020 1002.390 ;
        RECT 1714.020 1002.380 1717.020 1002.390 ;
        RECT 1894.020 1002.380 1897.020 1002.390 ;
        RECT 2074.020 1002.380 2077.020 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.300 1002.380 2934.300 1002.390 ;
        RECT -14.680 999.380 2934.300 1002.380 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 814.020 999.370 817.020 999.380 ;
        RECT 994.020 999.370 997.020 999.380 ;
        RECT 1174.020 999.370 1177.020 999.380 ;
        RECT 1354.020 999.370 1357.020 999.380 ;
        RECT 1534.020 999.370 1537.020 999.380 ;
        RECT 1714.020 999.370 1717.020 999.380 ;
        RECT 1894.020 999.370 1897.020 999.380 ;
        RECT 2074.020 999.370 2077.020 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.300 999.370 2934.300 999.380 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1534.020 822.380 1537.020 822.390 ;
        RECT 1714.020 822.380 1717.020 822.390 ;
        RECT 1894.020 822.380 1897.020 822.390 ;
        RECT 2074.020 822.380 2077.020 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.300 822.380 2934.300 822.390 ;
        RECT -14.680 819.380 2934.300 822.380 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1534.020 819.370 1537.020 819.380 ;
        RECT 1714.020 819.370 1717.020 819.380 ;
        RECT 1894.020 819.370 1897.020 819.380 ;
        RECT 2074.020 819.370 2077.020 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.300 819.370 2934.300 819.380 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1534.020 642.380 1537.020 642.390 ;
        RECT 1714.020 642.380 1717.020 642.390 ;
        RECT 1894.020 642.380 1897.020 642.390 ;
        RECT 2074.020 642.380 2077.020 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.300 642.380 2934.300 642.390 ;
        RECT -14.680 639.380 2934.300 642.380 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1534.020 639.370 1537.020 639.380 ;
        RECT 1714.020 639.370 1717.020 639.380 ;
        RECT 1894.020 639.370 1897.020 639.380 ;
        RECT 2074.020 639.370 2077.020 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.300 639.370 2934.300 639.380 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.300 462.380 2934.300 462.390 ;
        RECT -14.680 459.380 2934.300 462.380 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.300 459.370 2934.300 459.380 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.300 282.380 2934.300 282.390 ;
        RECT -14.680 279.380 2934.300 282.380 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.300 279.370 2934.300 279.380 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.300 102.380 2934.300 102.390 ;
        RECT -14.680 99.380 2934.300 102.380 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.300 99.370 2934.300 99.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT 22.020 -18.720 25.020 3538.400 ;
        RECT 202.020 -18.720 205.020 3538.400 ;
        RECT 382.020 -18.720 385.020 3538.400 ;
        RECT 562.020 -18.720 565.020 3538.400 ;
        RECT 742.020 -18.720 745.020 3538.400 ;
        RECT 922.020 -18.720 925.020 3538.400 ;
        RECT 1102.020 -18.720 1105.020 3538.400 ;
        RECT 1282.020 -18.720 1285.020 3538.400 ;
        RECT 1462.020 -18.720 1465.020 3538.400 ;
        RECT 1642.020 -18.720 1645.020 3538.400 ;
        RECT 1822.020 -18.720 1825.020 3538.400 ;
        RECT 2002.020 -18.720 2005.020 3538.400 ;
        RECT 2182.020 -18.720 2185.020 3538.400 ;
        RECT 2362.020 -18.720 2365.020 3538.400 ;
        RECT 2542.020 -18.720 2545.020 3538.400 ;
        RECT 2722.020 -18.720 2725.020 3538.400 ;
        RECT 2902.020 -18.720 2905.020 3538.400 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
      LAYER via4 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT -18.470 3449.090 -17.290 3450.270 ;
        RECT -18.470 3447.490 -17.290 3448.670 ;
        RECT -18.470 3269.090 -17.290 3270.270 ;
        RECT -18.470 3267.490 -17.290 3268.670 ;
        RECT -18.470 3089.090 -17.290 3090.270 ;
        RECT -18.470 3087.490 -17.290 3088.670 ;
        RECT -18.470 2909.090 -17.290 2910.270 ;
        RECT -18.470 2907.490 -17.290 2908.670 ;
        RECT -18.470 2729.090 -17.290 2730.270 ;
        RECT -18.470 2727.490 -17.290 2728.670 ;
        RECT -18.470 2549.090 -17.290 2550.270 ;
        RECT -18.470 2547.490 -17.290 2548.670 ;
        RECT -18.470 2369.090 -17.290 2370.270 ;
        RECT -18.470 2367.490 -17.290 2368.670 ;
        RECT -18.470 2189.090 -17.290 2190.270 ;
        RECT -18.470 2187.490 -17.290 2188.670 ;
        RECT -18.470 2009.090 -17.290 2010.270 ;
        RECT -18.470 2007.490 -17.290 2008.670 ;
        RECT -18.470 1829.090 -17.290 1830.270 ;
        RECT -18.470 1827.490 -17.290 1828.670 ;
        RECT -18.470 1649.090 -17.290 1650.270 ;
        RECT -18.470 1647.490 -17.290 1648.670 ;
        RECT -18.470 1469.090 -17.290 1470.270 ;
        RECT -18.470 1467.490 -17.290 1468.670 ;
        RECT -18.470 1289.090 -17.290 1290.270 ;
        RECT -18.470 1287.490 -17.290 1288.670 ;
        RECT -18.470 1109.090 -17.290 1110.270 ;
        RECT -18.470 1107.490 -17.290 1108.670 ;
        RECT -18.470 929.090 -17.290 930.270 ;
        RECT -18.470 927.490 -17.290 928.670 ;
        RECT -18.470 749.090 -17.290 750.270 ;
        RECT -18.470 747.490 -17.290 748.670 ;
        RECT -18.470 569.090 -17.290 570.270 ;
        RECT -18.470 567.490 -17.290 568.670 ;
        RECT -18.470 389.090 -17.290 390.270 ;
        RECT -18.470 387.490 -17.290 388.670 ;
        RECT -18.470 209.090 -17.290 210.270 ;
        RECT -18.470 207.490 -17.290 208.670 ;
        RECT -18.470 29.090 -17.290 30.270 ;
        RECT -18.470 27.490 -17.290 28.670 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 22.930 3532.410 24.110 3533.590 ;
        RECT 22.930 3530.810 24.110 3531.990 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.310 24.110 -11.130 ;
        RECT 22.930 -13.910 24.110 -12.730 ;
        RECT 202.930 3532.410 204.110 3533.590 ;
        RECT 202.930 3530.810 204.110 3531.990 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.310 204.110 -11.130 ;
        RECT 202.930 -13.910 204.110 -12.730 ;
        RECT 382.930 3532.410 384.110 3533.590 ;
        RECT 382.930 3530.810 384.110 3531.990 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 382.930 1829.090 384.110 1830.270 ;
        RECT 382.930 1827.490 384.110 1828.670 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.310 384.110 -11.130 ;
        RECT 382.930 -13.910 384.110 -12.730 ;
        RECT 562.930 3532.410 564.110 3533.590 ;
        RECT 562.930 3530.810 564.110 3531.990 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 562.930 2909.090 564.110 2910.270 ;
        RECT 562.930 2907.490 564.110 2908.670 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 562.930 2549.090 564.110 2550.270 ;
        RECT 562.930 2547.490 564.110 2548.670 ;
        RECT 562.930 2369.090 564.110 2370.270 ;
        RECT 562.930 2367.490 564.110 2368.670 ;
        RECT 562.930 2189.090 564.110 2190.270 ;
        RECT 562.930 2187.490 564.110 2188.670 ;
        RECT 562.930 2009.090 564.110 2010.270 ;
        RECT 562.930 2007.490 564.110 2008.670 ;
        RECT 562.930 1829.090 564.110 1830.270 ;
        RECT 562.930 1827.490 564.110 1828.670 ;
        RECT 562.930 1649.090 564.110 1650.270 ;
        RECT 562.930 1647.490 564.110 1648.670 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.310 564.110 -11.130 ;
        RECT 562.930 -13.910 564.110 -12.730 ;
        RECT 742.930 3532.410 744.110 3533.590 ;
        RECT 742.930 3530.810 744.110 3531.990 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 742.930 2549.090 744.110 2550.270 ;
        RECT 742.930 2547.490 744.110 2548.670 ;
        RECT 742.930 2369.090 744.110 2370.270 ;
        RECT 742.930 2367.490 744.110 2368.670 ;
        RECT 742.930 2189.090 744.110 2190.270 ;
        RECT 742.930 2187.490 744.110 2188.670 ;
        RECT 742.930 2009.090 744.110 2010.270 ;
        RECT 742.930 2007.490 744.110 2008.670 ;
        RECT 742.930 1829.090 744.110 1830.270 ;
        RECT 742.930 1827.490 744.110 1828.670 ;
        RECT 742.930 1649.090 744.110 1650.270 ;
        RECT 742.930 1647.490 744.110 1648.670 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.310 744.110 -11.130 ;
        RECT 742.930 -13.910 744.110 -12.730 ;
        RECT 922.930 3532.410 924.110 3533.590 ;
        RECT 922.930 3530.810 924.110 3531.990 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 922.930 2549.090 924.110 2550.270 ;
        RECT 922.930 2547.490 924.110 2548.670 ;
        RECT 922.930 2369.090 924.110 2370.270 ;
        RECT 922.930 2367.490 924.110 2368.670 ;
        RECT 922.930 2189.090 924.110 2190.270 ;
        RECT 922.930 2187.490 924.110 2188.670 ;
        RECT 922.930 2009.090 924.110 2010.270 ;
        RECT 922.930 2007.490 924.110 2008.670 ;
        RECT 922.930 1829.090 924.110 1830.270 ;
        RECT 922.930 1827.490 924.110 1828.670 ;
        RECT 922.930 1649.090 924.110 1650.270 ;
        RECT 922.930 1647.490 924.110 1648.670 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.310 924.110 -11.130 ;
        RECT 922.930 -13.910 924.110 -12.730 ;
        RECT 1102.930 3532.410 1104.110 3533.590 ;
        RECT 1102.930 3530.810 1104.110 3531.990 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1102.930 2909.090 1104.110 2910.270 ;
        RECT 1102.930 2907.490 1104.110 2908.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1102.930 2549.090 1104.110 2550.270 ;
        RECT 1102.930 2547.490 1104.110 2548.670 ;
        RECT 1102.930 2369.090 1104.110 2370.270 ;
        RECT 1102.930 2367.490 1104.110 2368.670 ;
        RECT 1102.930 2189.090 1104.110 2190.270 ;
        RECT 1102.930 2187.490 1104.110 2188.670 ;
        RECT 1102.930 2009.090 1104.110 2010.270 ;
        RECT 1102.930 2007.490 1104.110 2008.670 ;
        RECT 1102.930 1829.090 1104.110 1830.270 ;
        RECT 1102.930 1827.490 1104.110 1828.670 ;
        RECT 1102.930 1649.090 1104.110 1650.270 ;
        RECT 1102.930 1647.490 1104.110 1648.670 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.310 1104.110 -11.130 ;
        RECT 1102.930 -13.910 1104.110 -12.730 ;
        RECT 1282.930 3532.410 1284.110 3533.590 ;
        RECT 1282.930 3530.810 1284.110 3531.990 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1282.930 2909.090 1284.110 2910.270 ;
        RECT 1282.930 2907.490 1284.110 2908.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1282.930 2549.090 1284.110 2550.270 ;
        RECT 1282.930 2547.490 1284.110 2548.670 ;
        RECT 1282.930 2369.090 1284.110 2370.270 ;
        RECT 1282.930 2367.490 1284.110 2368.670 ;
        RECT 1282.930 2189.090 1284.110 2190.270 ;
        RECT 1282.930 2187.490 1284.110 2188.670 ;
        RECT 1282.930 2009.090 1284.110 2010.270 ;
        RECT 1282.930 2007.490 1284.110 2008.670 ;
        RECT 1282.930 1829.090 1284.110 1830.270 ;
        RECT 1282.930 1827.490 1284.110 1828.670 ;
        RECT 1282.930 1649.090 1284.110 1650.270 ;
        RECT 1282.930 1647.490 1284.110 1648.670 ;
        RECT 1282.930 1469.090 1284.110 1470.270 ;
        RECT 1282.930 1467.490 1284.110 1468.670 ;
        RECT 1282.930 1289.090 1284.110 1290.270 ;
        RECT 1282.930 1287.490 1284.110 1288.670 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.310 1284.110 -11.130 ;
        RECT 1282.930 -13.910 1284.110 -12.730 ;
        RECT 1462.930 3532.410 1464.110 3533.590 ;
        RECT 1462.930 3530.810 1464.110 3531.990 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 1462.930 2189.090 1464.110 2190.270 ;
        RECT 1462.930 2187.490 1464.110 2188.670 ;
        RECT 1462.930 2009.090 1464.110 2010.270 ;
        RECT 1462.930 2007.490 1464.110 2008.670 ;
        RECT 1462.930 1829.090 1464.110 1830.270 ;
        RECT 1462.930 1827.490 1464.110 1828.670 ;
        RECT 1462.930 1649.090 1464.110 1650.270 ;
        RECT 1462.930 1647.490 1464.110 1648.670 ;
        RECT 1462.930 1469.090 1464.110 1470.270 ;
        RECT 1462.930 1467.490 1464.110 1468.670 ;
        RECT 1462.930 1289.090 1464.110 1290.270 ;
        RECT 1462.930 1287.490 1464.110 1288.670 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.310 1464.110 -11.130 ;
        RECT 1462.930 -13.910 1464.110 -12.730 ;
        RECT 1642.930 3532.410 1644.110 3533.590 ;
        RECT 1642.930 3530.810 1644.110 3531.990 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1642.930 2909.090 1644.110 2910.270 ;
        RECT 1642.930 2907.490 1644.110 2908.670 ;
        RECT 1642.930 2729.090 1644.110 2730.270 ;
        RECT 1642.930 2727.490 1644.110 2728.670 ;
        RECT 1642.930 2549.090 1644.110 2550.270 ;
        RECT 1642.930 2547.490 1644.110 2548.670 ;
        RECT 1642.930 2369.090 1644.110 2370.270 ;
        RECT 1642.930 2367.490 1644.110 2368.670 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1642.930 2009.090 1644.110 2010.270 ;
        RECT 1642.930 2007.490 1644.110 2008.670 ;
        RECT 1642.930 1829.090 1644.110 1830.270 ;
        RECT 1642.930 1827.490 1644.110 1828.670 ;
        RECT 1642.930 1649.090 1644.110 1650.270 ;
        RECT 1642.930 1647.490 1644.110 1648.670 ;
        RECT 1642.930 1469.090 1644.110 1470.270 ;
        RECT 1642.930 1467.490 1644.110 1468.670 ;
        RECT 1642.930 1289.090 1644.110 1290.270 ;
        RECT 1642.930 1287.490 1644.110 1288.670 ;
        RECT 1642.930 1109.090 1644.110 1110.270 ;
        RECT 1642.930 1107.490 1644.110 1108.670 ;
        RECT 1642.930 929.090 1644.110 930.270 ;
        RECT 1642.930 927.490 1644.110 928.670 ;
        RECT 1642.930 749.090 1644.110 750.270 ;
        RECT 1642.930 747.490 1644.110 748.670 ;
        RECT 1642.930 569.090 1644.110 570.270 ;
        RECT 1642.930 567.490 1644.110 568.670 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.310 1644.110 -11.130 ;
        RECT 1642.930 -13.910 1644.110 -12.730 ;
        RECT 1822.930 3532.410 1824.110 3533.590 ;
        RECT 1822.930 3530.810 1824.110 3531.990 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 1822.930 2909.090 1824.110 2910.270 ;
        RECT 1822.930 2907.490 1824.110 2908.670 ;
        RECT 1822.930 2729.090 1824.110 2730.270 ;
        RECT 1822.930 2727.490 1824.110 2728.670 ;
        RECT 1822.930 2549.090 1824.110 2550.270 ;
        RECT 1822.930 2547.490 1824.110 2548.670 ;
        RECT 1822.930 2369.090 1824.110 2370.270 ;
        RECT 1822.930 2367.490 1824.110 2368.670 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1822.930 2009.090 1824.110 2010.270 ;
        RECT 1822.930 2007.490 1824.110 2008.670 ;
        RECT 1822.930 1829.090 1824.110 1830.270 ;
        RECT 1822.930 1827.490 1824.110 1828.670 ;
        RECT 1822.930 1649.090 1824.110 1650.270 ;
        RECT 1822.930 1647.490 1824.110 1648.670 ;
        RECT 1822.930 1469.090 1824.110 1470.270 ;
        RECT 1822.930 1467.490 1824.110 1468.670 ;
        RECT 1822.930 1289.090 1824.110 1290.270 ;
        RECT 1822.930 1287.490 1824.110 1288.670 ;
        RECT 1822.930 1109.090 1824.110 1110.270 ;
        RECT 1822.930 1107.490 1824.110 1108.670 ;
        RECT 1822.930 929.090 1824.110 930.270 ;
        RECT 1822.930 927.490 1824.110 928.670 ;
        RECT 1822.930 749.090 1824.110 750.270 ;
        RECT 1822.930 747.490 1824.110 748.670 ;
        RECT 1822.930 569.090 1824.110 570.270 ;
        RECT 1822.930 567.490 1824.110 568.670 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.310 1824.110 -11.130 ;
        RECT 1822.930 -13.910 1824.110 -12.730 ;
        RECT 2002.930 3532.410 2004.110 3533.590 ;
        RECT 2002.930 3530.810 2004.110 3531.990 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 2002.930 2369.090 2004.110 2370.270 ;
        RECT 2002.930 2367.490 2004.110 2368.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 2002.930 2009.090 2004.110 2010.270 ;
        RECT 2002.930 2007.490 2004.110 2008.670 ;
        RECT 2002.930 1829.090 2004.110 1830.270 ;
        RECT 2002.930 1827.490 2004.110 1828.670 ;
        RECT 2002.930 1649.090 2004.110 1650.270 ;
        RECT 2002.930 1647.490 2004.110 1648.670 ;
        RECT 2002.930 1469.090 2004.110 1470.270 ;
        RECT 2002.930 1467.490 2004.110 1468.670 ;
        RECT 2002.930 1289.090 2004.110 1290.270 ;
        RECT 2002.930 1287.490 2004.110 1288.670 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 2002.930 929.090 2004.110 930.270 ;
        RECT 2002.930 927.490 2004.110 928.670 ;
        RECT 2002.930 749.090 2004.110 750.270 ;
        RECT 2002.930 747.490 2004.110 748.670 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.310 2004.110 -11.130 ;
        RECT 2002.930 -13.910 2004.110 -12.730 ;
        RECT 2182.930 3532.410 2184.110 3533.590 ;
        RECT 2182.930 3530.810 2184.110 3531.990 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2182.930 2909.090 2184.110 2910.270 ;
        RECT 2182.930 2907.490 2184.110 2908.670 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2182.930 2369.090 2184.110 2370.270 ;
        RECT 2182.930 2367.490 2184.110 2368.670 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2182.930 2009.090 2184.110 2010.270 ;
        RECT 2182.930 2007.490 2184.110 2008.670 ;
        RECT 2182.930 1829.090 2184.110 1830.270 ;
        RECT 2182.930 1827.490 2184.110 1828.670 ;
        RECT 2182.930 1649.090 2184.110 1650.270 ;
        RECT 2182.930 1647.490 2184.110 1648.670 ;
        RECT 2182.930 1469.090 2184.110 1470.270 ;
        RECT 2182.930 1467.490 2184.110 1468.670 ;
        RECT 2182.930 1289.090 2184.110 1290.270 ;
        RECT 2182.930 1287.490 2184.110 1288.670 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 2182.930 929.090 2184.110 930.270 ;
        RECT 2182.930 927.490 2184.110 928.670 ;
        RECT 2182.930 749.090 2184.110 750.270 ;
        RECT 2182.930 747.490 2184.110 748.670 ;
        RECT 2182.930 569.090 2184.110 570.270 ;
        RECT 2182.930 567.490 2184.110 568.670 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.310 2184.110 -11.130 ;
        RECT 2182.930 -13.910 2184.110 -12.730 ;
        RECT 2362.930 3532.410 2364.110 3533.590 ;
        RECT 2362.930 3530.810 2364.110 3531.990 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2362.930 2909.090 2364.110 2910.270 ;
        RECT 2362.930 2907.490 2364.110 2908.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2362.930 2009.090 2364.110 2010.270 ;
        RECT 2362.930 2007.490 2364.110 2008.670 ;
        RECT 2362.930 1829.090 2364.110 1830.270 ;
        RECT 2362.930 1827.490 2364.110 1828.670 ;
        RECT 2362.930 1649.090 2364.110 1650.270 ;
        RECT 2362.930 1647.490 2364.110 1648.670 ;
        RECT 2362.930 1469.090 2364.110 1470.270 ;
        RECT 2362.930 1467.490 2364.110 1468.670 ;
        RECT 2362.930 1289.090 2364.110 1290.270 ;
        RECT 2362.930 1287.490 2364.110 1288.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2362.930 929.090 2364.110 930.270 ;
        RECT 2362.930 927.490 2364.110 928.670 ;
        RECT 2362.930 749.090 2364.110 750.270 ;
        RECT 2362.930 747.490 2364.110 748.670 ;
        RECT 2362.930 569.090 2364.110 570.270 ;
        RECT 2362.930 567.490 2364.110 568.670 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.310 2364.110 -11.130 ;
        RECT 2362.930 -13.910 2364.110 -12.730 ;
        RECT 2542.930 3532.410 2544.110 3533.590 ;
        RECT 2542.930 3530.810 2544.110 3531.990 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.310 2544.110 -11.130 ;
        RECT 2542.930 -13.910 2544.110 -12.730 ;
        RECT 2722.930 3532.410 2724.110 3533.590 ;
        RECT 2722.930 3530.810 2724.110 3531.990 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.310 2724.110 -11.130 ;
        RECT 2722.930 -13.910 2724.110 -12.730 ;
        RECT 2902.930 3532.410 2904.110 3533.590 ;
        RECT 2902.930 3530.810 2904.110 3531.990 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.310 2904.110 -11.130 ;
        RECT 2902.930 -13.910 2904.110 -12.730 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2936.910 3449.090 2938.090 3450.270 ;
        RECT 2936.910 3447.490 2938.090 3448.670 ;
        RECT 2936.910 3269.090 2938.090 3270.270 ;
        RECT 2936.910 3267.490 2938.090 3268.670 ;
        RECT 2936.910 3089.090 2938.090 3090.270 ;
        RECT 2936.910 3087.490 2938.090 3088.670 ;
        RECT 2936.910 2909.090 2938.090 2910.270 ;
        RECT 2936.910 2907.490 2938.090 2908.670 ;
        RECT 2936.910 2729.090 2938.090 2730.270 ;
        RECT 2936.910 2727.490 2938.090 2728.670 ;
        RECT 2936.910 2549.090 2938.090 2550.270 ;
        RECT 2936.910 2547.490 2938.090 2548.670 ;
        RECT 2936.910 2369.090 2938.090 2370.270 ;
        RECT 2936.910 2367.490 2938.090 2368.670 ;
        RECT 2936.910 2189.090 2938.090 2190.270 ;
        RECT 2936.910 2187.490 2938.090 2188.670 ;
        RECT 2936.910 2009.090 2938.090 2010.270 ;
        RECT 2936.910 2007.490 2938.090 2008.670 ;
        RECT 2936.910 1829.090 2938.090 1830.270 ;
        RECT 2936.910 1827.490 2938.090 1828.670 ;
        RECT 2936.910 1649.090 2938.090 1650.270 ;
        RECT 2936.910 1647.490 2938.090 1648.670 ;
        RECT 2936.910 1469.090 2938.090 1470.270 ;
        RECT 2936.910 1467.490 2938.090 1468.670 ;
        RECT 2936.910 1289.090 2938.090 1290.270 ;
        RECT 2936.910 1287.490 2938.090 1288.670 ;
        RECT 2936.910 1109.090 2938.090 1110.270 ;
        RECT 2936.910 1107.490 2938.090 1108.670 ;
        RECT 2936.910 929.090 2938.090 930.270 ;
        RECT 2936.910 927.490 2938.090 928.670 ;
        RECT 2936.910 749.090 2938.090 750.270 ;
        RECT 2936.910 747.490 2938.090 748.670 ;
        RECT 2936.910 569.090 2938.090 570.270 ;
        RECT 2936.910 567.490 2938.090 568.670 ;
        RECT 2936.910 389.090 2938.090 390.270 ;
        RECT 2936.910 387.490 2938.090 388.670 ;
        RECT 2936.910 209.090 2938.090 210.270 ;
        RECT 2936.910 207.490 2938.090 208.670 ;
        RECT 2936.910 29.090 2938.090 30.270 ;
        RECT 2936.910 27.490 2938.090 28.670 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
      LAYER met5 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 22.020 3533.700 25.020 3533.710 ;
        RECT 202.020 3533.700 205.020 3533.710 ;
        RECT 382.020 3533.700 385.020 3533.710 ;
        RECT 562.020 3533.700 565.020 3533.710 ;
        RECT 742.020 3533.700 745.020 3533.710 ;
        RECT 922.020 3533.700 925.020 3533.710 ;
        RECT 1102.020 3533.700 1105.020 3533.710 ;
        RECT 1282.020 3533.700 1285.020 3533.710 ;
        RECT 1462.020 3533.700 1465.020 3533.710 ;
        RECT 1642.020 3533.700 1645.020 3533.710 ;
        RECT 1822.020 3533.700 1825.020 3533.710 ;
        RECT 2002.020 3533.700 2005.020 3533.710 ;
        RECT 2182.020 3533.700 2185.020 3533.710 ;
        RECT 2362.020 3533.700 2365.020 3533.710 ;
        RECT 2542.020 3533.700 2545.020 3533.710 ;
        RECT 2722.020 3533.700 2725.020 3533.710 ;
        RECT 2902.020 3533.700 2905.020 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 22.020 3530.690 25.020 3530.700 ;
        RECT 202.020 3530.690 205.020 3530.700 ;
        RECT 382.020 3530.690 385.020 3530.700 ;
        RECT 562.020 3530.690 565.020 3530.700 ;
        RECT 742.020 3530.690 745.020 3530.700 ;
        RECT 922.020 3530.690 925.020 3530.700 ;
        RECT 1102.020 3530.690 1105.020 3530.700 ;
        RECT 1282.020 3530.690 1285.020 3530.700 ;
        RECT 1462.020 3530.690 1465.020 3530.700 ;
        RECT 1642.020 3530.690 1645.020 3530.700 ;
        RECT 1822.020 3530.690 1825.020 3530.700 ;
        RECT 2002.020 3530.690 2005.020 3530.700 ;
        RECT 2182.020 3530.690 2185.020 3530.700 ;
        RECT 2362.020 3530.690 2365.020 3530.700 ;
        RECT 2542.020 3530.690 2545.020 3530.700 ;
        RECT 2722.020 3530.690 2725.020 3530.700 ;
        RECT 2902.020 3530.690 2905.020 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -19.380 3450.380 -16.380 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2936.000 3450.380 2939.000 3450.390 ;
        RECT -24.080 3447.380 2943.700 3450.380 ;
        RECT -19.380 3447.370 -16.380 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2936.000 3447.370 2939.000 3447.380 ;
        RECT -19.380 3270.380 -16.380 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2936.000 3270.380 2939.000 3270.390 ;
        RECT -24.080 3267.380 2943.700 3270.380 ;
        RECT -19.380 3267.370 -16.380 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2936.000 3267.370 2939.000 3267.380 ;
        RECT -19.380 3090.380 -16.380 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2936.000 3090.380 2939.000 3090.390 ;
        RECT -24.080 3087.380 2943.700 3090.380 ;
        RECT -19.380 3087.370 -16.380 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2936.000 3087.370 2939.000 3087.380 ;
        RECT -19.380 2910.380 -16.380 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 562.020 2910.380 565.020 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1102.020 2910.380 1105.020 2910.390 ;
        RECT 1282.020 2910.380 1285.020 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1642.020 2910.380 1645.020 2910.390 ;
        RECT 1822.020 2910.380 1825.020 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2182.020 2910.380 2185.020 2910.390 ;
        RECT 2362.020 2910.380 2365.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2936.000 2910.380 2939.000 2910.390 ;
        RECT -24.080 2907.380 2943.700 2910.380 ;
        RECT -19.380 2907.370 -16.380 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 562.020 2907.370 565.020 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1102.020 2907.370 1105.020 2907.380 ;
        RECT 1282.020 2907.370 1285.020 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1642.020 2907.370 1645.020 2907.380 ;
        RECT 1822.020 2907.370 1825.020 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2182.020 2907.370 2185.020 2907.380 ;
        RECT 2362.020 2907.370 2365.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2936.000 2907.370 2939.000 2907.380 ;
        RECT -19.380 2730.380 -16.380 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 1642.020 2730.380 1645.020 2730.390 ;
        RECT 1822.020 2730.380 1825.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2936.000 2730.380 2939.000 2730.390 ;
        RECT -24.080 2727.380 2943.700 2730.380 ;
        RECT -19.380 2727.370 -16.380 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 1642.020 2727.370 1645.020 2727.380 ;
        RECT 1822.020 2727.370 1825.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2936.000 2727.370 2939.000 2727.380 ;
        RECT -19.380 2550.380 -16.380 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 562.020 2550.380 565.020 2550.390 ;
        RECT 742.020 2550.380 745.020 2550.390 ;
        RECT 922.020 2550.380 925.020 2550.390 ;
        RECT 1102.020 2550.380 1105.020 2550.390 ;
        RECT 1282.020 2550.380 1285.020 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 1642.020 2550.380 1645.020 2550.390 ;
        RECT 1822.020 2550.380 1825.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2936.000 2550.380 2939.000 2550.390 ;
        RECT -24.080 2547.380 2943.700 2550.380 ;
        RECT -19.380 2547.370 -16.380 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 562.020 2547.370 565.020 2547.380 ;
        RECT 742.020 2547.370 745.020 2547.380 ;
        RECT 922.020 2547.370 925.020 2547.380 ;
        RECT 1102.020 2547.370 1105.020 2547.380 ;
        RECT 1282.020 2547.370 1285.020 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 1642.020 2547.370 1645.020 2547.380 ;
        RECT 1822.020 2547.370 1825.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2936.000 2547.370 2939.000 2547.380 ;
        RECT -19.380 2370.380 -16.380 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 562.020 2370.380 565.020 2370.390 ;
        RECT 742.020 2370.380 745.020 2370.390 ;
        RECT 922.020 2370.380 925.020 2370.390 ;
        RECT 1102.020 2370.380 1105.020 2370.390 ;
        RECT 1282.020 2370.380 1285.020 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 1642.020 2370.380 1645.020 2370.390 ;
        RECT 1822.020 2370.380 1825.020 2370.390 ;
        RECT 2002.020 2370.380 2005.020 2370.390 ;
        RECT 2182.020 2370.380 2185.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2936.000 2370.380 2939.000 2370.390 ;
        RECT -24.080 2367.380 2943.700 2370.380 ;
        RECT -19.380 2367.370 -16.380 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 562.020 2367.370 565.020 2367.380 ;
        RECT 742.020 2367.370 745.020 2367.380 ;
        RECT 922.020 2367.370 925.020 2367.380 ;
        RECT 1102.020 2367.370 1105.020 2367.380 ;
        RECT 1282.020 2367.370 1285.020 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 1642.020 2367.370 1645.020 2367.380 ;
        RECT 1822.020 2367.370 1825.020 2367.380 ;
        RECT 2002.020 2367.370 2005.020 2367.380 ;
        RECT 2182.020 2367.370 2185.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2936.000 2367.370 2939.000 2367.380 ;
        RECT -19.380 2190.380 -16.380 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 562.020 2190.380 565.020 2190.390 ;
        RECT 742.020 2190.380 745.020 2190.390 ;
        RECT 922.020 2190.380 925.020 2190.390 ;
        RECT 1102.020 2190.380 1105.020 2190.390 ;
        RECT 1282.020 2190.380 1285.020 2190.390 ;
        RECT 1462.020 2190.380 1465.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2936.000 2190.380 2939.000 2190.390 ;
        RECT -24.080 2187.380 2943.700 2190.380 ;
        RECT -19.380 2187.370 -16.380 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 562.020 2187.370 565.020 2187.380 ;
        RECT 742.020 2187.370 745.020 2187.380 ;
        RECT 922.020 2187.370 925.020 2187.380 ;
        RECT 1102.020 2187.370 1105.020 2187.380 ;
        RECT 1282.020 2187.370 1285.020 2187.380 ;
        RECT 1462.020 2187.370 1465.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2936.000 2187.370 2939.000 2187.380 ;
        RECT -19.380 2010.380 -16.380 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 562.020 2010.380 565.020 2010.390 ;
        RECT 742.020 2010.380 745.020 2010.390 ;
        RECT 922.020 2010.380 925.020 2010.390 ;
        RECT 1102.020 2010.380 1105.020 2010.390 ;
        RECT 1282.020 2010.380 1285.020 2010.390 ;
        RECT 1462.020 2010.380 1465.020 2010.390 ;
        RECT 1642.020 2010.380 1645.020 2010.390 ;
        RECT 1822.020 2010.380 1825.020 2010.390 ;
        RECT 2002.020 2010.380 2005.020 2010.390 ;
        RECT 2182.020 2010.380 2185.020 2010.390 ;
        RECT 2362.020 2010.380 2365.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2936.000 2010.380 2939.000 2010.390 ;
        RECT -24.080 2007.380 2943.700 2010.380 ;
        RECT -19.380 2007.370 -16.380 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 562.020 2007.370 565.020 2007.380 ;
        RECT 742.020 2007.370 745.020 2007.380 ;
        RECT 922.020 2007.370 925.020 2007.380 ;
        RECT 1102.020 2007.370 1105.020 2007.380 ;
        RECT 1282.020 2007.370 1285.020 2007.380 ;
        RECT 1462.020 2007.370 1465.020 2007.380 ;
        RECT 1642.020 2007.370 1645.020 2007.380 ;
        RECT 1822.020 2007.370 1825.020 2007.380 ;
        RECT 2002.020 2007.370 2005.020 2007.380 ;
        RECT 2182.020 2007.370 2185.020 2007.380 ;
        RECT 2362.020 2007.370 2365.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2936.000 2007.370 2939.000 2007.380 ;
        RECT -19.380 1830.380 -16.380 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 382.020 1830.380 385.020 1830.390 ;
        RECT 562.020 1830.380 565.020 1830.390 ;
        RECT 742.020 1830.380 745.020 1830.390 ;
        RECT 922.020 1830.380 925.020 1830.390 ;
        RECT 1102.020 1830.380 1105.020 1830.390 ;
        RECT 1282.020 1830.380 1285.020 1830.390 ;
        RECT 1462.020 1830.380 1465.020 1830.390 ;
        RECT 1642.020 1830.380 1645.020 1830.390 ;
        RECT 1822.020 1830.380 1825.020 1830.390 ;
        RECT 2002.020 1830.380 2005.020 1830.390 ;
        RECT 2182.020 1830.380 2185.020 1830.390 ;
        RECT 2362.020 1830.380 2365.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2936.000 1830.380 2939.000 1830.390 ;
        RECT -24.080 1827.380 2943.700 1830.380 ;
        RECT -19.380 1827.370 -16.380 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 382.020 1827.370 385.020 1827.380 ;
        RECT 562.020 1827.370 565.020 1827.380 ;
        RECT 742.020 1827.370 745.020 1827.380 ;
        RECT 922.020 1827.370 925.020 1827.380 ;
        RECT 1102.020 1827.370 1105.020 1827.380 ;
        RECT 1282.020 1827.370 1285.020 1827.380 ;
        RECT 1462.020 1827.370 1465.020 1827.380 ;
        RECT 1642.020 1827.370 1645.020 1827.380 ;
        RECT 1822.020 1827.370 1825.020 1827.380 ;
        RECT 2002.020 1827.370 2005.020 1827.380 ;
        RECT 2182.020 1827.370 2185.020 1827.380 ;
        RECT 2362.020 1827.370 2365.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2936.000 1827.370 2939.000 1827.380 ;
        RECT -19.380 1650.380 -16.380 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 562.020 1650.380 565.020 1650.390 ;
        RECT 742.020 1650.380 745.020 1650.390 ;
        RECT 922.020 1650.380 925.020 1650.390 ;
        RECT 1102.020 1650.380 1105.020 1650.390 ;
        RECT 1282.020 1650.380 1285.020 1650.390 ;
        RECT 1462.020 1650.380 1465.020 1650.390 ;
        RECT 1642.020 1650.380 1645.020 1650.390 ;
        RECT 1822.020 1650.380 1825.020 1650.390 ;
        RECT 2002.020 1650.380 2005.020 1650.390 ;
        RECT 2182.020 1650.380 2185.020 1650.390 ;
        RECT 2362.020 1650.380 2365.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2936.000 1650.380 2939.000 1650.390 ;
        RECT -24.080 1647.380 2943.700 1650.380 ;
        RECT -19.380 1647.370 -16.380 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 562.020 1647.370 565.020 1647.380 ;
        RECT 742.020 1647.370 745.020 1647.380 ;
        RECT 922.020 1647.370 925.020 1647.380 ;
        RECT 1102.020 1647.370 1105.020 1647.380 ;
        RECT 1282.020 1647.370 1285.020 1647.380 ;
        RECT 1462.020 1647.370 1465.020 1647.380 ;
        RECT 1642.020 1647.370 1645.020 1647.380 ;
        RECT 1822.020 1647.370 1825.020 1647.380 ;
        RECT 2002.020 1647.370 2005.020 1647.380 ;
        RECT 2182.020 1647.370 2185.020 1647.380 ;
        RECT 2362.020 1647.370 2365.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2936.000 1647.370 2939.000 1647.380 ;
        RECT -19.380 1470.380 -16.380 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 1282.020 1470.380 1285.020 1470.390 ;
        RECT 1462.020 1470.380 1465.020 1470.390 ;
        RECT 1642.020 1470.380 1645.020 1470.390 ;
        RECT 1822.020 1470.380 1825.020 1470.390 ;
        RECT 2002.020 1470.380 2005.020 1470.390 ;
        RECT 2182.020 1470.380 2185.020 1470.390 ;
        RECT 2362.020 1470.380 2365.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2936.000 1470.380 2939.000 1470.390 ;
        RECT -24.080 1467.380 2943.700 1470.380 ;
        RECT -19.380 1467.370 -16.380 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 1282.020 1467.370 1285.020 1467.380 ;
        RECT 1462.020 1467.370 1465.020 1467.380 ;
        RECT 1642.020 1467.370 1645.020 1467.380 ;
        RECT 1822.020 1467.370 1825.020 1467.380 ;
        RECT 2002.020 1467.370 2005.020 1467.380 ;
        RECT 2182.020 1467.370 2185.020 1467.380 ;
        RECT 2362.020 1467.370 2365.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2936.000 1467.370 2939.000 1467.380 ;
        RECT -19.380 1290.380 -16.380 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 1282.020 1290.380 1285.020 1290.390 ;
        RECT 1462.020 1290.380 1465.020 1290.390 ;
        RECT 1642.020 1290.380 1645.020 1290.390 ;
        RECT 1822.020 1290.380 1825.020 1290.390 ;
        RECT 2002.020 1290.380 2005.020 1290.390 ;
        RECT 2182.020 1290.380 2185.020 1290.390 ;
        RECT 2362.020 1290.380 2365.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2936.000 1290.380 2939.000 1290.390 ;
        RECT -24.080 1287.380 2943.700 1290.380 ;
        RECT -19.380 1287.370 -16.380 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 1282.020 1287.370 1285.020 1287.380 ;
        RECT 1462.020 1287.370 1465.020 1287.380 ;
        RECT 1642.020 1287.370 1645.020 1287.380 ;
        RECT 1822.020 1287.370 1825.020 1287.380 ;
        RECT 2002.020 1287.370 2005.020 1287.380 ;
        RECT 2182.020 1287.370 2185.020 1287.380 ;
        RECT 2362.020 1287.370 2365.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2936.000 1287.370 2939.000 1287.380 ;
        RECT -19.380 1110.380 -16.380 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1642.020 1110.380 1645.020 1110.390 ;
        RECT 1822.020 1110.380 1825.020 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2936.000 1110.380 2939.000 1110.390 ;
        RECT -24.080 1107.380 2943.700 1110.380 ;
        RECT -19.380 1107.370 -16.380 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1642.020 1107.370 1645.020 1107.380 ;
        RECT 1822.020 1107.370 1825.020 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2936.000 1107.370 2939.000 1107.380 ;
        RECT -19.380 930.380 -16.380 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 1642.020 930.380 1645.020 930.390 ;
        RECT 1822.020 930.380 1825.020 930.390 ;
        RECT 2002.020 930.380 2005.020 930.390 ;
        RECT 2182.020 930.380 2185.020 930.390 ;
        RECT 2362.020 930.380 2365.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2936.000 930.380 2939.000 930.390 ;
        RECT -24.080 927.380 2943.700 930.380 ;
        RECT -19.380 927.370 -16.380 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 1642.020 927.370 1645.020 927.380 ;
        RECT 1822.020 927.370 1825.020 927.380 ;
        RECT 2002.020 927.370 2005.020 927.380 ;
        RECT 2182.020 927.370 2185.020 927.380 ;
        RECT 2362.020 927.370 2365.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2936.000 927.370 2939.000 927.380 ;
        RECT -19.380 750.380 -16.380 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 1642.020 750.380 1645.020 750.390 ;
        RECT 1822.020 750.380 1825.020 750.390 ;
        RECT 2002.020 750.380 2005.020 750.390 ;
        RECT 2182.020 750.380 2185.020 750.390 ;
        RECT 2362.020 750.380 2365.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2936.000 750.380 2939.000 750.390 ;
        RECT -24.080 747.380 2943.700 750.380 ;
        RECT -19.380 747.370 -16.380 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 1642.020 747.370 1645.020 747.380 ;
        RECT 1822.020 747.370 1825.020 747.380 ;
        RECT 2002.020 747.370 2005.020 747.380 ;
        RECT 2182.020 747.370 2185.020 747.380 ;
        RECT 2362.020 747.370 2365.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2936.000 747.370 2939.000 747.380 ;
        RECT -19.380 570.380 -16.380 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1642.020 570.380 1645.020 570.390 ;
        RECT 1822.020 570.380 1825.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2182.020 570.380 2185.020 570.390 ;
        RECT 2362.020 570.380 2365.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2936.000 570.380 2939.000 570.390 ;
        RECT -24.080 567.380 2943.700 570.380 ;
        RECT -19.380 567.370 -16.380 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1642.020 567.370 1645.020 567.380 ;
        RECT 1822.020 567.370 1825.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2182.020 567.370 2185.020 567.380 ;
        RECT 2362.020 567.370 2365.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2936.000 567.370 2939.000 567.380 ;
        RECT -19.380 390.380 -16.380 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2936.000 390.380 2939.000 390.390 ;
        RECT -24.080 387.380 2943.700 390.380 ;
        RECT -19.380 387.370 -16.380 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2936.000 387.370 2939.000 387.380 ;
        RECT -19.380 210.380 -16.380 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2936.000 210.380 2939.000 210.390 ;
        RECT -24.080 207.380 2943.700 210.380 ;
        RECT -19.380 207.370 -16.380 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2936.000 207.370 2939.000 207.380 ;
        RECT -19.380 30.380 -16.380 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2936.000 30.380 2939.000 30.390 ;
        RECT -24.080 27.380 2943.700 30.380 ;
        RECT -19.380 27.370 -16.380 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2936.000 27.370 2939.000 27.380 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 22.020 -11.020 25.020 -11.010 ;
        RECT 202.020 -11.020 205.020 -11.010 ;
        RECT 382.020 -11.020 385.020 -11.010 ;
        RECT 562.020 -11.020 565.020 -11.010 ;
        RECT 742.020 -11.020 745.020 -11.010 ;
        RECT 922.020 -11.020 925.020 -11.010 ;
        RECT 1102.020 -11.020 1105.020 -11.010 ;
        RECT 1282.020 -11.020 1285.020 -11.010 ;
        RECT 1462.020 -11.020 1465.020 -11.010 ;
        RECT 1642.020 -11.020 1645.020 -11.010 ;
        RECT 1822.020 -11.020 1825.020 -11.010 ;
        RECT 2002.020 -11.020 2005.020 -11.010 ;
        RECT 2182.020 -11.020 2185.020 -11.010 ;
        RECT 2362.020 -11.020 2365.020 -11.010 ;
        RECT 2542.020 -11.020 2545.020 -11.010 ;
        RECT 2722.020 -11.020 2725.020 -11.010 ;
        RECT 2902.020 -11.020 2905.020 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 22.020 -14.030 25.020 -14.020 ;
        RECT 202.020 -14.030 205.020 -14.020 ;
        RECT 382.020 -14.030 385.020 -14.020 ;
        RECT 562.020 -14.030 565.020 -14.020 ;
        RECT 742.020 -14.030 745.020 -14.020 ;
        RECT 922.020 -14.030 925.020 -14.020 ;
        RECT 1102.020 -14.030 1105.020 -14.020 ;
        RECT 1282.020 -14.030 1285.020 -14.020 ;
        RECT 1462.020 -14.030 1465.020 -14.020 ;
        RECT 1642.020 -14.030 1645.020 -14.020 ;
        RECT 1822.020 -14.030 1825.020 -14.020 ;
        RECT 2002.020 -14.030 2005.020 -14.020 ;
        RECT 2182.020 -14.030 2185.020 -14.020 ;
        RECT 2362.020 -14.030 2365.020 -14.020 ;
        RECT 2542.020 -14.030 2545.020 -14.020 ;
        RECT 2722.020 -14.030 2725.020 -14.020 ;
        RECT 2902.020 -14.030 2905.020 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT 112.020 -18.720 115.020 3538.400 ;
        RECT 292.020 -18.720 295.020 3538.400 ;
        RECT 472.020 -18.720 475.020 3538.400 ;
        RECT 652.020 -18.720 655.020 3538.400 ;
        RECT 832.020 -18.720 835.020 3538.400 ;
        RECT 1012.020 -18.720 1015.020 3538.400 ;
        RECT 1192.020 -18.720 1195.020 3538.400 ;
        RECT 1372.020 -18.720 1375.020 3538.400 ;
        RECT 1552.020 -18.720 1555.020 3538.400 ;
        RECT 1732.020 -18.720 1735.020 3538.400 ;
        RECT 1912.020 -18.720 1915.020 3538.400 ;
        RECT 2092.020 -18.720 2095.020 3538.400 ;
        RECT 2272.020 -18.720 2275.020 3538.400 ;
        RECT 2452.020 -18.720 2455.020 3538.400 ;
        RECT 2632.020 -18.720 2635.020 3538.400 ;
        RECT 2812.020 -18.720 2815.020 3538.400 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
      LAYER via4 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT -23.170 3359.090 -21.990 3360.270 ;
        RECT -23.170 3357.490 -21.990 3358.670 ;
        RECT -23.170 3179.090 -21.990 3180.270 ;
        RECT -23.170 3177.490 -21.990 3178.670 ;
        RECT -23.170 2999.090 -21.990 3000.270 ;
        RECT -23.170 2997.490 -21.990 2998.670 ;
        RECT -23.170 2819.090 -21.990 2820.270 ;
        RECT -23.170 2817.490 -21.990 2818.670 ;
        RECT -23.170 2639.090 -21.990 2640.270 ;
        RECT -23.170 2637.490 -21.990 2638.670 ;
        RECT -23.170 2459.090 -21.990 2460.270 ;
        RECT -23.170 2457.490 -21.990 2458.670 ;
        RECT -23.170 2279.090 -21.990 2280.270 ;
        RECT -23.170 2277.490 -21.990 2278.670 ;
        RECT -23.170 2099.090 -21.990 2100.270 ;
        RECT -23.170 2097.490 -21.990 2098.670 ;
        RECT -23.170 1919.090 -21.990 1920.270 ;
        RECT -23.170 1917.490 -21.990 1918.670 ;
        RECT -23.170 1739.090 -21.990 1740.270 ;
        RECT -23.170 1737.490 -21.990 1738.670 ;
        RECT -23.170 1559.090 -21.990 1560.270 ;
        RECT -23.170 1557.490 -21.990 1558.670 ;
        RECT -23.170 1379.090 -21.990 1380.270 ;
        RECT -23.170 1377.490 -21.990 1378.670 ;
        RECT -23.170 1199.090 -21.990 1200.270 ;
        RECT -23.170 1197.490 -21.990 1198.670 ;
        RECT -23.170 1019.090 -21.990 1020.270 ;
        RECT -23.170 1017.490 -21.990 1018.670 ;
        RECT -23.170 839.090 -21.990 840.270 ;
        RECT -23.170 837.490 -21.990 838.670 ;
        RECT -23.170 659.090 -21.990 660.270 ;
        RECT -23.170 657.490 -21.990 658.670 ;
        RECT -23.170 479.090 -21.990 480.270 ;
        RECT -23.170 477.490 -21.990 478.670 ;
        RECT -23.170 299.090 -21.990 300.270 ;
        RECT -23.170 297.490 -21.990 298.670 ;
        RECT -23.170 119.090 -21.990 120.270 ;
        RECT -23.170 117.490 -21.990 118.670 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 112.930 3537.110 114.110 3538.290 ;
        RECT 112.930 3535.510 114.110 3536.690 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -17.010 114.110 -15.830 ;
        RECT 112.930 -18.610 114.110 -17.430 ;
        RECT 292.930 3537.110 294.110 3538.290 ;
        RECT 292.930 3535.510 294.110 3536.690 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -17.010 294.110 -15.830 ;
        RECT 292.930 -18.610 294.110 -17.430 ;
        RECT 472.930 3537.110 474.110 3538.290 ;
        RECT 472.930 3535.510 474.110 3536.690 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 472.930 2999.090 474.110 3000.270 ;
        RECT 472.930 2997.490 474.110 2998.670 ;
        RECT 472.930 2819.090 474.110 2820.270 ;
        RECT 472.930 2817.490 474.110 2818.670 ;
        RECT 472.930 2639.090 474.110 2640.270 ;
        RECT 472.930 2637.490 474.110 2638.670 ;
        RECT 472.930 2459.090 474.110 2460.270 ;
        RECT 472.930 2457.490 474.110 2458.670 ;
        RECT 472.930 2279.090 474.110 2280.270 ;
        RECT 472.930 2277.490 474.110 2278.670 ;
        RECT 472.930 2099.090 474.110 2100.270 ;
        RECT 472.930 2097.490 474.110 2098.670 ;
        RECT 472.930 1919.090 474.110 1920.270 ;
        RECT 472.930 1917.490 474.110 1918.670 ;
        RECT 472.930 1739.090 474.110 1740.270 ;
        RECT 472.930 1737.490 474.110 1738.670 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -17.010 474.110 -15.830 ;
        RECT 472.930 -18.610 474.110 -17.430 ;
        RECT 652.930 3537.110 654.110 3538.290 ;
        RECT 652.930 3535.510 654.110 3536.690 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 652.930 2999.090 654.110 3000.270 ;
        RECT 652.930 2997.490 654.110 2998.670 ;
        RECT 652.930 2819.090 654.110 2820.270 ;
        RECT 652.930 2817.490 654.110 2818.670 ;
        RECT 652.930 2639.090 654.110 2640.270 ;
        RECT 652.930 2637.490 654.110 2638.670 ;
        RECT 652.930 2459.090 654.110 2460.270 ;
        RECT 652.930 2457.490 654.110 2458.670 ;
        RECT 652.930 2279.090 654.110 2280.270 ;
        RECT 652.930 2277.490 654.110 2278.670 ;
        RECT 652.930 2099.090 654.110 2100.270 ;
        RECT 652.930 2097.490 654.110 2098.670 ;
        RECT 652.930 1919.090 654.110 1920.270 ;
        RECT 652.930 1917.490 654.110 1918.670 ;
        RECT 652.930 1739.090 654.110 1740.270 ;
        RECT 652.930 1737.490 654.110 1738.670 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -17.010 654.110 -15.830 ;
        RECT 652.930 -18.610 654.110 -17.430 ;
        RECT 832.930 3537.110 834.110 3538.290 ;
        RECT 832.930 3535.510 834.110 3536.690 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 832.930 2639.090 834.110 2640.270 ;
        RECT 832.930 2637.490 834.110 2638.670 ;
        RECT 832.930 2459.090 834.110 2460.270 ;
        RECT 832.930 2457.490 834.110 2458.670 ;
        RECT 832.930 2279.090 834.110 2280.270 ;
        RECT 832.930 2277.490 834.110 2278.670 ;
        RECT 832.930 2099.090 834.110 2100.270 ;
        RECT 832.930 2097.490 834.110 2098.670 ;
        RECT 832.930 1919.090 834.110 1920.270 ;
        RECT 832.930 1917.490 834.110 1918.670 ;
        RECT 832.930 1739.090 834.110 1740.270 ;
        RECT 832.930 1737.490 834.110 1738.670 ;
        RECT 832.930 1559.090 834.110 1560.270 ;
        RECT 832.930 1557.490 834.110 1558.670 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -17.010 834.110 -15.830 ;
        RECT 832.930 -18.610 834.110 -17.430 ;
        RECT 1012.930 3537.110 1014.110 3538.290 ;
        RECT 1012.930 3535.510 1014.110 3536.690 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1012.930 2999.090 1014.110 3000.270 ;
        RECT 1012.930 2997.490 1014.110 2998.670 ;
        RECT 1012.930 2819.090 1014.110 2820.270 ;
        RECT 1012.930 2817.490 1014.110 2818.670 ;
        RECT 1012.930 2639.090 1014.110 2640.270 ;
        RECT 1012.930 2637.490 1014.110 2638.670 ;
        RECT 1012.930 2459.090 1014.110 2460.270 ;
        RECT 1012.930 2457.490 1014.110 2458.670 ;
        RECT 1012.930 2279.090 1014.110 2280.270 ;
        RECT 1012.930 2277.490 1014.110 2278.670 ;
        RECT 1012.930 2099.090 1014.110 2100.270 ;
        RECT 1012.930 2097.490 1014.110 2098.670 ;
        RECT 1012.930 1919.090 1014.110 1920.270 ;
        RECT 1012.930 1917.490 1014.110 1918.670 ;
        RECT 1012.930 1739.090 1014.110 1740.270 ;
        RECT 1012.930 1737.490 1014.110 1738.670 ;
        RECT 1012.930 1559.090 1014.110 1560.270 ;
        RECT 1012.930 1557.490 1014.110 1558.670 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -17.010 1014.110 -15.830 ;
        RECT 1012.930 -18.610 1014.110 -17.430 ;
        RECT 1192.930 3537.110 1194.110 3538.290 ;
        RECT 1192.930 3535.510 1194.110 3536.690 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1192.930 2999.090 1194.110 3000.270 ;
        RECT 1192.930 2997.490 1194.110 2998.670 ;
        RECT 1192.930 2819.090 1194.110 2820.270 ;
        RECT 1192.930 2817.490 1194.110 2818.670 ;
        RECT 1192.930 2639.090 1194.110 2640.270 ;
        RECT 1192.930 2637.490 1194.110 2638.670 ;
        RECT 1192.930 2459.090 1194.110 2460.270 ;
        RECT 1192.930 2457.490 1194.110 2458.670 ;
        RECT 1192.930 2279.090 1194.110 2280.270 ;
        RECT 1192.930 2277.490 1194.110 2278.670 ;
        RECT 1192.930 2099.090 1194.110 2100.270 ;
        RECT 1192.930 2097.490 1194.110 2098.670 ;
        RECT 1192.930 1919.090 1194.110 1920.270 ;
        RECT 1192.930 1917.490 1194.110 1918.670 ;
        RECT 1192.930 1739.090 1194.110 1740.270 ;
        RECT 1192.930 1737.490 1194.110 1738.670 ;
        RECT 1192.930 1559.090 1194.110 1560.270 ;
        RECT 1192.930 1557.490 1194.110 1558.670 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -17.010 1194.110 -15.830 ;
        RECT 1192.930 -18.610 1194.110 -17.430 ;
        RECT 1372.930 3537.110 1374.110 3538.290 ;
        RECT 1372.930 3535.510 1374.110 3536.690 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1372.930 2639.090 1374.110 2640.270 ;
        RECT 1372.930 2637.490 1374.110 2638.670 ;
        RECT 1372.930 2459.090 1374.110 2460.270 ;
        RECT 1372.930 2457.490 1374.110 2458.670 ;
        RECT 1372.930 2279.090 1374.110 2280.270 ;
        RECT 1372.930 2277.490 1374.110 2278.670 ;
        RECT 1372.930 2099.090 1374.110 2100.270 ;
        RECT 1372.930 2097.490 1374.110 2098.670 ;
        RECT 1372.930 1919.090 1374.110 1920.270 ;
        RECT 1372.930 1917.490 1374.110 1918.670 ;
        RECT 1372.930 1739.090 1374.110 1740.270 ;
        RECT 1372.930 1737.490 1374.110 1738.670 ;
        RECT 1372.930 1559.090 1374.110 1560.270 ;
        RECT 1372.930 1557.490 1374.110 1558.670 ;
        RECT 1372.930 1379.090 1374.110 1380.270 ;
        RECT 1372.930 1377.490 1374.110 1378.670 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -17.010 1374.110 -15.830 ;
        RECT 1372.930 -18.610 1374.110 -17.430 ;
        RECT 1552.930 3537.110 1554.110 3538.290 ;
        RECT 1552.930 3535.510 1554.110 3536.690 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1552.930 2999.090 1554.110 3000.270 ;
        RECT 1552.930 2997.490 1554.110 2998.670 ;
        RECT 1552.930 2819.090 1554.110 2820.270 ;
        RECT 1552.930 2817.490 1554.110 2818.670 ;
        RECT 1552.930 2639.090 1554.110 2640.270 ;
        RECT 1552.930 2637.490 1554.110 2638.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 1552.930 2099.090 1554.110 2100.270 ;
        RECT 1552.930 2097.490 1554.110 2098.670 ;
        RECT 1552.930 1919.090 1554.110 1920.270 ;
        RECT 1552.930 1917.490 1554.110 1918.670 ;
        RECT 1552.930 1739.090 1554.110 1740.270 ;
        RECT 1552.930 1737.490 1554.110 1738.670 ;
        RECT 1552.930 1559.090 1554.110 1560.270 ;
        RECT 1552.930 1557.490 1554.110 1558.670 ;
        RECT 1552.930 1379.090 1554.110 1380.270 ;
        RECT 1552.930 1377.490 1554.110 1378.670 ;
        RECT 1552.930 1199.090 1554.110 1200.270 ;
        RECT 1552.930 1197.490 1554.110 1198.670 ;
        RECT 1552.930 1019.090 1554.110 1020.270 ;
        RECT 1552.930 1017.490 1554.110 1018.670 ;
        RECT 1552.930 839.090 1554.110 840.270 ;
        RECT 1552.930 837.490 1554.110 838.670 ;
        RECT 1552.930 659.090 1554.110 660.270 ;
        RECT 1552.930 657.490 1554.110 658.670 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -17.010 1554.110 -15.830 ;
        RECT 1552.930 -18.610 1554.110 -17.430 ;
        RECT 1732.930 3537.110 1734.110 3538.290 ;
        RECT 1732.930 3535.510 1734.110 3536.690 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1732.930 2999.090 1734.110 3000.270 ;
        RECT 1732.930 2997.490 1734.110 2998.670 ;
        RECT 1732.930 2819.090 1734.110 2820.270 ;
        RECT 1732.930 2817.490 1734.110 2818.670 ;
        RECT 1732.930 2639.090 1734.110 2640.270 ;
        RECT 1732.930 2637.490 1734.110 2638.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 1732.930 2279.090 1734.110 2280.270 ;
        RECT 1732.930 2277.490 1734.110 2278.670 ;
        RECT 1732.930 2099.090 1734.110 2100.270 ;
        RECT 1732.930 2097.490 1734.110 2098.670 ;
        RECT 1732.930 1919.090 1734.110 1920.270 ;
        RECT 1732.930 1917.490 1734.110 1918.670 ;
        RECT 1732.930 1739.090 1734.110 1740.270 ;
        RECT 1732.930 1737.490 1734.110 1738.670 ;
        RECT 1732.930 1559.090 1734.110 1560.270 ;
        RECT 1732.930 1557.490 1734.110 1558.670 ;
        RECT 1732.930 1379.090 1734.110 1380.270 ;
        RECT 1732.930 1377.490 1734.110 1378.670 ;
        RECT 1732.930 1199.090 1734.110 1200.270 ;
        RECT 1732.930 1197.490 1734.110 1198.670 ;
        RECT 1732.930 1019.090 1734.110 1020.270 ;
        RECT 1732.930 1017.490 1734.110 1018.670 ;
        RECT 1732.930 839.090 1734.110 840.270 ;
        RECT 1732.930 837.490 1734.110 838.670 ;
        RECT 1732.930 659.090 1734.110 660.270 ;
        RECT 1732.930 657.490 1734.110 658.670 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -17.010 1734.110 -15.830 ;
        RECT 1732.930 -18.610 1734.110 -17.430 ;
        RECT 1912.930 3537.110 1914.110 3538.290 ;
        RECT 1912.930 3535.510 1914.110 3536.690 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 1912.930 2999.090 1914.110 3000.270 ;
        RECT 1912.930 2997.490 1914.110 2998.670 ;
        RECT 1912.930 2819.090 1914.110 2820.270 ;
        RECT 1912.930 2817.490 1914.110 2818.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 1912.930 2279.090 1914.110 2280.270 ;
        RECT 1912.930 2277.490 1914.110 2278.670 ;
        RECT 1912.930 2099.090 1914.110 2100.270 ;
        RECT 1912.930 2097.490 1914.110 2098.670 ;
        RECT 1912.930 1919.090 1914.110 1920.270 ;
        RECT 1912.930 1917.490 1914.110 1918.670 ;
        RECT 1912.930 1739.090 1914.110 1740.270 ;
        RECT 1912.930 1737.490 1914.110 1738.670 ;
        RECT 1912.930 1559.090 1914.110 1560.270 ;
        RECT 1912.930 1557.490 1914.110 1558.670 ;
        RECT 1912.930 1379.090 1914.110 1380.270 ;
        RECT 1912.930 1377.490 1914.110 1378.670 ;
        RECT 1912.930 1199.090 1914.110 1200.270 ;
        RECT 1912.930 1197.490 1914.110 1198.670 ;
        RECT 1912.930 1019.090 1914.110 1020.270 ;
        RECT 1912.930 1017.490 1914.110 1018.670 ;
        RECT 1912.930 839.090 1914.110 840.270 ;
        RECT 1912.930 837.490 1914.110 838.670 ;
        RECT 1912.930 659.090 1914.110 660.270 ;
        RECT 1912.930 657.490 1914.110 658.670 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -17.010 1914.110 -15.830 ;
        RECT 1912.930 -18.610 1914.110 -17.430 ;
        RECT 2092.930 3537.110 2094.110 3538.290 ;
        RECT 2092.930 3535.510 2094.110 3536.690 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 2092.930 1919.090 2094.110 1920.270 ;
        RECT 2092.930 1917.490 2094.110 1918.670 ;
        RECT 2092.930 1739.090 2094.110 1740.270 ;
        RECT 2092.930 1737.490 2094.110 1738.670 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2092.930 1379.090 2094.110 1380.270 ;
        RECT 2092.930 1377.490 2094.110 1378.670 ;
        RECT 2092.930 1199.090 2094.110 1200.270 ;
        RECT 2092.930 1197.490 2094.110 1198.670 ;
        RECT 2092.930 1019.090 2094.110 1020.270 ;
        RECT 2092.930 1017.490 2094.110 1018.670 ;
        RECT 2092.930 839.090 2094.110 840.270 ;
        RECT 2092.930 837.490 2094.110 838.670 ;
        RECT 2092.930 659.090 2094.110 660.270 ;
        RECT 2092.930 657.490 2094.110 658.670 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -17.010 2094.110 -15.830 ;
        RECT 2092.930 -18.610 2094.110 -17.430 ;
        RECT 2272.930 3537.110 2274.110 3538.290 ;
        RECT 2272.930 3535.510 2274.110 3536.690 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2272.930 2999.090 2274.110 3000.270 ;
        RECT 2272.930 2997.490 2274.110 2998.670 ;
        RECT 2272.930 2819.090 2274.110 2820.270 ;
        RECT 2272.930 2817.490 2274.110 2818.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2272.930 1919.090 2274.110 1920.270 ;
        RECT 2272.930 1917.490 2274.110 1918.670 ;
        RECT 2272.930 1739.090 2274.110 1740.270 ;
        RECT 2272.930 1737.490 2274.110 1738.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2272.930 1379.090 2274.110 1380.270 ;
        RECT 2272.930 1377.490 2274.110 1378.670 ;
        RECT 2272.930 1199.090 2274.110 1200.270 ;
        RECT 2272.930 1197.490 2274.110 1198.670 ;
        RECT 2272.930 1019.090 2274.110 1020.270 ;
        RECT 2272.930 1017.490 2274.110 1018.670 ;
        RECT 2272.930 839.090 2274.110 840.270 ;
        RECT 2272.930 837.490 2274.110 838.670 ;
        RECT 2272.930 659.090 2274.110 660.270 ;
        RECT 2272.930 657.490 2274.110 658.670 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -17.010 2274.110 -15.830 ;
        RECT 2272.930 -18.610 2274.110 -17.430 ;
        RECT 2452.930 3537.110 2454.110 3538.290 ;
        RECT 2452.930 3535.510 2454.110 3536.690 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2452.930 2999.090 2454.110 3000.270 ;
        RECT 2452.930 2997.490 2454.110 2998.670 ;
        RECT 2452.930 2819.090 2454.110 2820.270 ;
        RECT 2452.930 2817.490 2454.110 2818.670 ;
        RECT 2452.930 2639.090 2454.110 2640.270 ;
        RECT 2452.930 2637.490 2454.110 2638.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2452.930 1919.090 2454.110 1920.270 ;
        RECT 2452.930 1917.490 2454.110 1918.670 ;
        RECT 2452.930 1739.090 2454.110 1740.270 ;
        RECT 2452.930 1737.490 2454.110 1738.670 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2452.930 1379.090 2454.110 1380.270 ;
        RECT 2452.930 1377.490 2454.110 1378.670 ;
        RECT 2452.930 1199.090 2454.110 1200.270 ;
        RECT 2452.930 1197.490 2454.110 1198.670 ;
        RECT 2452.930 1019.090 2454.110 1020.270 ;
        RECT 2452.930 1017.490 2454.110 1018.670 ;
        RECT 2452.930 839.090 2454.110 840.270 ;
        RECT 2452.930 837.490 2454.110 838.670 ;
        RECT 2452.930 659.090 2454.110 660.270 ;
        RECT 2452.930 657.490 2454.110 658.670 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -17.010 2454.110 -15.830 ;
        RECT 2452.930 -18.610 2454.110 -17.430 ;
        RECT 2632.930 3537.110 2634.110 3538.290 ;
        RECT 2632.930 3535.510 2634.110 3536.690 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -17.010 2634.110 -15.830 ;
        RECT 2632.930 -18.610 2634.110 -17.430 ;
        RECT 2812.930 3537.110 2814.110 3538.290 ;
        RECT 2812.930 3535.510 2814.110 3536.690 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -17.010 2814.110 -15.830 ;
        RECT 2812.930 -18.610 2814.110 -17.430 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT 2941.610 3359.090 2942.790 3360.270 ;
        RECT 2941.610 3357.490 2942.790 3358.670 ;
        RECT 2941.610 3179.090 2942.790 3180.270 ;
        RECT 2941.610 3177.490 2942.790 3178.670 ;
        RECT 2941.610 2999.090 2942.790 3000.270 ;
        RECT 2941.610 2997.490 2942.790 2998.670 ;
        RECT 2941.610 2819.090 2942.790 2820.270 ;
        RECT 2941.610 2817.490 2942.790 2818.670 ;
        RECT 2941.610 2639.090 2942.790 2640.270 ;
        RECT 2941.610 2637.490 2942.790 2638.670 ;
        RECT 2941.610 2459.090 2942.790 2460.270 ;
        RECT 2941.610 2457.490 2942.790 2458.670 ;
        RECT 2941.610 2279.090 2942.790 2280.270 ;
        RECT 2941.610 2277.490 2942.790 2278.670 ;
        RECT 2941.610 2099.090 2942.790 2100.270 ;
        RECT 2941.610 2097.490 2942.790 2098.670 ;
        RECT 2941.610 1919.090 2942.790 1920.270 ;
        RECT 2941.610 1917.490 2942.790 1918.670 ;
        RECT 2941.610 1739.090 2942.790 1740.270 ;
        RECT 2941.610 1737.490 2942.790 1738.670 ;
        RECT 2941.610 1559.090 2942.790 1560.270 ;
        RECT 2941.610 1557.490 2942.790 1558.670 ;
        RECT 2941.610 1379.090 2942.790 1380.270 ;
        RECT 2941.610 1377.490 2942.790 1378.670 ;
        RECT 2941.610 1199.090 2942.790 1200.270 ;
        RECT 2941.610 1197.490 2942.790 1198.670 ;
        RECT 2941.610 1019.090 2942.790 1020.270 ;
        RECT 2941.610 1017.490 2942.790 1018.670 ;
        RECT 2941.610 839.090 2942.790 840.270 ;
        RECT 2941.610 837.490 2942.790 838.670 ;
        RECT 2941.610 659.090 2942.790 660.270 ;
        RECT 2941.610 657.490 2942.790 658.670 ;
        RECT 2941.610 479.090 2942.790 480.270 ;
        RECT 2941.610 477.490 2942.790 478.670 ;
        RECT 2941.610 299.090 2942.790 300.270 ;
        RECT 2941.610 297.490 2942.790 298.670 ;
        RECT 2941.610 119.090 2942.790 120.270 ;
        RECT 2941.610 117.490 2942.790 118.670 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
      LAYER met5 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 112.020 3538.400 115.020 3538.410 ;
        RECT 292.020 3538.400 295.020 3538.410 ;
        RECT 472.020 3538.400 475.020 3538.410 ;
        RECT 652.020 3538.400 655.020 3538.410 ;
        RECT 832.020 3538.400 835.020 3538.410 ;
        RECT 1012.020 3538.400 1015.020 3538.410 ;
        RECT 1192.020 3538.400 1195.020 3538.410 ;
        RECT 1372.020 3538.400 1375.020 3538.410 ;
        RECT 1552.020 3538.400 1555.020 3538.410 ;
        RECT 1732.020 3538.400 1735.020 3538.410 ;
        RECT 1912.020 3538.400 1915.020 3538.410 ;
        RECT 2092.020 3538.400 2095.020 3538.410 ;
        RECT 2272.020 3538.400 2275.020 3538.410 ;
        RECT 2452.020 3538.400 2455.020 3538.410 ;
        RECT 2632.020 3538.400 2635.020 3538.410 ;
        RECT 2812.020 3538.400 2815.020 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 112.020 3535.390 115.020 3535.400 ;
        RECT 292.020 3535.390 295.020 3535.400 ;
        RECT 472.020 3535.390 475.020 3535.400 ;
        RECT 652.020 3535.390 655.020 3535.400 ;
        RECT 832.020 3535.390 835.020 3535.400 ;
        RECT 1012.020 3535.390 1015.020 3535.400 ;
        RECT 1192.020 3535.390 1195.020 3535.400 ;
        RECT 1372.020 3535.390 1375.020 3535.400 ;
        RECT 1552.020 3535.390 1555.020 3535.400 ;
        RECT 1732.020 3535.390 1735.020 3535.400 ;
        RECT 1912.020 3535.390 1915.020 3535.400 ;
        RECT 2092.020 3535.390 2095.020 3535.400 ;
        RECT 2272.020 3535.390 2275.020 3535.400 ;
        RECT 2452.020 3535.390 2455.020 3535.400 ;
        RECT 2632.020 3535.390 2635.020 3535.400 ;
        RECT 2812.020 3535.390 2815.020 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -24.080 3360.380 -21.080 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.700 3360.380 2943.700 3360.390 ;
        RECT -24.080 3357.380 2943.700 3360.380 ;
        RECT -24.080 3357.370 -21.080 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.700 3357.370 2943.700 3357.380 ;
        RECT -24.080 3180.380 -21.080 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.700 3180.380 2943.700 3180.390 ;
        RECT -24.080 3177.380 2943.700 3180.380 ;
        RECT -24.080 3177.370 -21.080 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.700 3177.370 2943.700 3177.380 ;
        RECT -24.080 3000.380 -21.080 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 472.020 3000.380 475.020 3000.390 ;
        RECT 652.020 3000.380 655.020 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1012.020 3000.380 1015.020 3000.390 ;
        RECT 1192.020 3000.380 1195.020 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1552.020 3000.380 1555.020 3000.390 ;
        RECT 1732.020 3000.380 1735.020 3000.390 ;
        RECT 1912.020 3000.380 1915.020 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2272.020 3000.380 2275.020 3000.390 ;
        RECT 2452.020 3000.380 2455.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.700 3000.380 2943.700 3000.390 ;
        RECT -24.080 2997.380 2943.700 3000.380 ;
        RECT -24.080 2997.370 -21.080 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 472.020 2997.370 475.020 2997.380 ;
        RECT 652.020 2997.370 655.020 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1012.020 2997.370 1015.020 2997.380 ;
        RECT 1192.020 2997.370 1195.020 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1552.020 2997.370 1555.020 2997.380 ;
        RECT 1732.020 2997.370 1735.020 2997.380 ;
        RECT 1912.020 2997.370 1915.020 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2272.020 2997.370 2275.020 2997.380 ;
        RECT 2452.020 2997.370 2455.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.700 2997.370 2943.700 2997.380 ;
        RECT -24.080 2820.380 -21.080 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 472.020 2820.380 475.020 2820.390 ;
        RECT 652.020 2820.380 655.020 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1012.020 2820.380 1015.020 2820.390 ;
        RECT 1192.020 2820.380 1195.020 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1552.020 2820.380 1555.020 2820.390 ;
        RECT 1732.020 2820.380 1735.020 2820.390 ;
        RECT 1912.020 2820.380 1915.020 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2272.020 2820.380 2275.020 2820.390 ;
        RECT 2452.020 2820.380 2455.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.700 2820.380 2943.700 2820.390 ;
        RECT -24.080 2817.380 2943.700 2820.380 ;
        RECT -24.080 2817.370 -21.080 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 472.020 2817.370 475.020 2817.380 ;
        RECT 652.020 2817.370 655.020 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1012.020 2817.370 1015.020 2817.380 ;
        RECT 1192.020 2817.370 1195.020 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1552.020 2817.370 1555.020 2817.380 ;
        RECT 1732.020 2817.370 1735.020 2817.380 ;
        RECT 1912.020 2817.370 1915.020 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2272.020 2817.370 2275.020 2817.380 ;
        RECT 2452.020 2817.370 2455.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.700 2817.370 2943.700 2817.380 ;
        RECT -24.080 2640.380 -21.080 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 472.020 2640.380 475.020 2640.390 ;
        RECT 652.020 2640.380 655.020 2640.390 ;
        RECT 832.020 2640.380 835.020 2640.390 ;
        RECT 1012.020 2640.380 1015.020 2640.390 ;
        RECT 1192.020 2640.380 1195.020 2640.390 ;
        RECT 1372.020 2640.380 1375.020 2640.390 ;
        RECT 1552.020 2640.380 1555.020 2640.390 ;
        RECT 1732.020 2640.380 1735.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2452.020 2640.380 2455.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.700 2640.380 2943.700 2640.390 ;
        RECT -24.080 2637.380 2943.700 2640.380 ;
        RECT -24.080 2637.370 -21.080 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 472.020 2637.370 475.020 2637.380 ;
        RECT 652.020 2637.370 655.020 2637.380 ;
        RECT 832.020 2637.370 835.020 2637.380 ;
        RECT 1012.020 2637.370 1015.020 2637.380 ;
        RECT 1192.020 2637.370 1195.020 2637.380 ;
        RECT 1372.020 2637.370 1375.020 2637.380 ;
        RECT 1552.020 2637.370 1555.020 2637.380 ;
        RECT 1732.020 2637.370 1735.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2452.020 2637.370 2455.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.700 2637.370 2943.700 2637.380 ;
        RECT -24.080 2460.380 -21.080 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 472.020 2460.380 475.020 2460.390 ;
        RECT 652.020 2460.380 655.020 2460.390 ;
        RECT 832.020 2460.380 835.020 2460.390 ;
        RECT 1012.020 2460.380 1015.020 2460.390 ;
        RECT 1192.020 2460.380 1195.020 2460.390 ;
        RECT 1372.020 2460.380 1375.020 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.700 2460.380 2943.700 2460.390 ;
        RECT -24.080 2457.380 2943.700 2460.380 ;
        RECT -24.080 2457.370 -21.080 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 472.020 2457.370 475.020 2457.380 ;
        RECT 652.020 2457.370 655.020 2457.380 ;
        RECT 832.020 2457.370 835.020 2457.380 ;
        RECT 1012.020 2457.370 1015.020 2457.380 ;
        RECT 1192.020 2457.370 1195.020 2457.380 ;
        RECT 1372.020 2457.370 1375.020 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.700 2457.370 2943.700 2457.380 ;
        RECT -24.080 2280.380 -21.080 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 472.020 2280.380 475.020 2280.390 ;
        RECT 652.020 2280.380 655.020 2280.390 ;
        RECT 832.020 2280.380 835.020 2280.390 ;
        RECT 1012.020 2280.380 1015.020 2280.390 ;
        RECT 1192.020 2280.380 1195.020 2280.390 ;
        RECT 1372.020 2280.380 1375.020 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 1732.020 2280.380 1735.020 2280.390 ;
        RECT 1912.020 2280.380 1915.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.700 2280.380 2943.700 2280.390 ;
        RECT -24.080 2277.380 2943.700 2280.380 ;
        RECT -24.080 2277.370 -21.080 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 472.020 2277.370 475.020 2277.380 ;
        RECT 652.020 2277.370 655.020 2277.380 ;
        RECT 832.020 2277.370 835.020 2277.380 ;
        RECT 1012.020 2277.370 1015.020 2277.380 ;
        RECT 1192.020 2277.370 1195.020 2277.380 ;
        RECT 1372.020 2277.370 1375.020 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 1732.020 2277.370 1735.020 2277.380 ;
        RECT 1912.020 2277.370 1915.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.700 2277.370 2943.700 2277.380 ;
        RECT -24.080 2100.380 -21.080 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 472.020 2100.380 475.020 2100.390 ;
        RECT 652.020 2100.380 655.020 2100.390 ;
        RECT 832.020 2100.380 835.020 2100.390 ;
        RECT 1012.020 2100.380 1015.020 2100.390 ;
        RECT 1192.020 2100.380 1195.020 2100.390 ;
        RECT 1372.020 2100.380 1375.020 2100.390 ;
        RECT 1552.020 2100.380 1555.020 2100.390 ;
        RECT 1732.020 2100.380 1735.020 2100.390 ;
        RECT 1912.020 2100.380 1915.020 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.700 2100.380 2943.700 2100.390 ;
        RECT -24.080 2097.380 2943.700 2100.380 ;
        RECT -24.080 2097.370 -21.080 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 472.020 2097.370 475.020 2097.380 ;
        RECT 652.020 2097.370 655.020 2097.380 ;
        RECT 832.020 2097.370 835.020 2097.380 ;
        RECT 1012.020 2097.370 1015.020 2097.380 ;
        RECT 1192.020 2097.370 1195.020 2097.380 ;
        RECT 1372.020 2097.370 1375.020 2097.380 ;
        RECT 1552.020 2097.370 1555.020 2097.380 ;
        RECT 1732.020 2097.370 1735.020 2097.380 ;
        RECT 1912.020 2097.370 1915.020 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.700 2097.370 2943.700 2097.380 ;
        RECT -24.080 1920.380 -21.080 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 472.020 1920.380 475.020 1920.390 ;
        RECT 652.020 1920.380 655.020 1920.390 ;
        RECT 832.020 1920.380 835.020 1920.390 ;
        RECT 1012.020 1920.380 1015.020 1920.390 ;
        RECT 1192.020 1920.380 1195.020 1920.390 ;
        RECT 1372.020 1920.380 1375.020 1920.390 ;
        RECT 1552.020 1920.380 1555.020 1920.390 ;
        RECT 1732.020 1920.380 1735.020 1920.390 ;
        RECT 1912.020 1920.380 1915.020 1920.390 ;
        RECT 2092.020 1920.380 2095.020 1920.390 ;
        RECT 2272.020 1920.380 2275.020 1920.390 ;
        RECT 2452.020 1920.380 2455.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.700 1920.380 2943.700 1920.390 ;
        RECT -24.080 1917.380 2943.700 1920.380 ;
        RECT -24.080 1917.370 -21.080 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 472.020 1917.370 475.020 1917.380 ;
        RECT 652.020 1917.370 655.020 1917.380 ;
        RECT 832.020 1917.370 835.020 1917.380 ;
        RECT 1012.020 1917.370 1015.020 1917.380 ;
        RECT 1192.020 1917.370 1195.020 1917.380 ;
        RECT 1372.020 1917.370 1375.020 1917.380 ;
        RECT 1552.020 1917.370 1555.020 1917.380 ;
        RECT 1732.020 1917.370 1735.020 1917.380 ;
        RECT 1912.020 1917.370 1915.020 1917.380 ;
        RECT 2092.020 1917.370 2095.020 1917.380 ;
        RECT 2272.020 1917.370 2275.020 1917.380 ;
        RECT 2452.020 1917.370 2455.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.700 1917.370 2943.700 1917.380 ;
        RECT -24.080 1740.380 -21.080 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 472.020 1740.380 475.020 1740.390 ;
        RECT 652.020 1740.380 655.020 1740.390 ;
        RECT 832.020 1740.380 835.020 1740.390 ;
        RECT 1012.020 1740.380 1015.020 1740.390 ;
        RECT 1192.020 1740.380 1195.020 1740.390 ;
        RECT 1372.020 1740.380 1375.020 1740.390 ;
        RECT 1552.020 1740.380 1555.020 1740.390 ;
        RECT 1732.020 1740.380 1735.020 1740.390 ;
        RECT 1912.020 1740.380 1915.020 1740.390 ;
        RECT 2092.020 1740.380 2095.020 1740.390 ;
        RECT 2272.020 1740.380 2275.020 1740.390 ;
        RECT 2452.020 1740.380 2455.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.700 1740.380 2943.700 1740.390 ;
        RECT -24.080 1737.380 2943.700 1740.380 ;
        RECT -24.080 1737.370 -21.080 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 472.020 1737.370 475.020 1737.380 ;
        RECT 652.020 1737.370 655.020 1737.380 ;
        RECT 832.020 1737.370 835.020 1737.380 ;
        RECT 1012.020 1737.370 1015.020 1737.380 ;
        RECT 1192.020 1737.370 1195.020 1737.380 ;
        RECT 1372.020 1737.370 1375.020 1737.380 ;
        RECT 1552.020 1737.370 1555.020 1737.380 ;
        RECT 1732.020 1737.370 1735.020 1737.380 ;
        RECT 1912.020 1737.370 1915.020 1737.380 ;
        RECT 2092.020 1737.370 2095.020 1737.380 ;
        RECT 2272.020 1737.370 2275.020 1737.380 ;
        RECT 2452.020 1737.370 2455.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.700 1737.370 2943.700 1737.380 ;
        RECT -24.080 1560.380 -21.080 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 832.020 1560.380 835.020 1560.390 ;
        RECT 1012.020 1560.380 1015.020 1560.390 ;
        RECT 1192.020 1560.380 1195.020 1560.390 ;
        RECT 1372.020 1560.380 1375.020 1560.390 ;
        RECT 1552.020 1560.380 1555.020 1560.390 ;
        RECT 1732.020 1560.380 1735.020 1560.390 ;
        RECT 1912.020 1560.380 1915.020 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.700 1560.380 2943.700 1560.390 ;
        RECT -24.080 1557.380 2943.700 1560.380 ;
        RECT -24.080 1557.370 -21.080 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 832.020 1557.370 835.020 1557.380 ;
        RECT 1012.020 1557.370 1015.020 1557.380 ;
        RECT 1192.020 1557.370 1195.020 1557.380 ;
        RECT 1372.020 1557.370 1375.020 1557.380 ;
        RECT 1552.020 1557.370 1555.020 1557.380 ;
        RECT 1732.020 1557.370 1735.020 1557.380 ;
        RECT 1912.020 1557.370 1915.020 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.700 1557.370 2943.700 1557.380 ;
        RECT -24.080 1380.380 -21.080 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 1372.020 1380.380 1375.020 1380.390 ;
        RECT 1552.020 1380.380 1555.020 1380.390 ;
        RECT 1732.020 1380.380 1735.020 1380.390 ;
        RECT 1912.020 1380.380 1915.020 1380.390 ;
        RECT 2092.020 1380.380 2095.020 1380.390 ;
        RECT 2272.020 1380.380 2275.020 1380.390 ;
        RECT 2452.020 1380.380 2455.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.700 1380.380 2943.700 1380.390 ;
        RECT -24.080 1377.380 2943.700 1380.380 ;
        RECT -24.080 1377.370 -21.080 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 1372.020 1377.370 1375.020 1377.380 ;
        RECT 1552.020 1377.370 1555.020 1377.380 ;
        RECT 1732.020 1377.370 1735.020 1377.380 ;
        RECT 1912.020 1377.370 1915.020 1377.380 ;
        RECT 2092.020 1377.370 2095.020 1377.380 ;
        RECT 2272.020 1377.370 2275.020 1377.380 ;
        RECT 2452.020 1377.370 2455.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.700 1377.370 2943.700 1377.380 ;
        RECT -24.080 1200.380 -21.080 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 1552.020 1200.380 1555.020 1200.390 ;
        RECT 1732.020 1200.380 1735.020 1200.390 ;
        RECT 1912.020 1200.380 1915.020 1200.390 ;
        RECT 2092.020 1200.380 2095.020 1200.390 ;
        RECT 2272.020 1200.380 2275.020 1200.390 ;
        RECT 2452.020 1200.380 2455.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.700 1200.380 2943.700 1200.390 ;
        RECT -24.080 1197.380 2943.700 1200.380 ;
        RECT -24.080 1197.370 -21.080 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 1552.020 1197.370 1555.020 1197.380 ;
        RECT 1732.020 1197.370 1735.020 1197.380 ;
        RECT 1912.020 1197.370 1915.020 1197.380 ;
        RECT 2092.020 1197.370 2095.020 1197.380 ;
        RECT 2272.020 1197.370 2275.020 1197.380 ;
        RECT 2452.020 1197.370 2455.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.700 1197.370 2943.700 1197.380 ;
        RECT -24.080 1020.380 -21.080 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1552.020 1020.380 1555.020 1020.390 ;
        RECT 1732.020 1020.380 1735.020 1020.390 ;
        RECT 1912.020 1020.380 1915.020 1020.390 ;
        RECT 2092.020 1020.380 2095.020 1020.390 ;
        RECT 2272.020 1020.380 2275.020 1020.390 ;
        RECT 2452.020 1020.380 2455.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.700 1020.380 2943.700 1020.390 ;
        RECT -24.080 1017.380 2943.700 1020.380 ;
        RECT -24.080 1017.370 -21.080 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1552.020 1017.370 1555.020 1017.380 ;
        RECT 1732.020 1017.370 1735.020 1017.380 ;
        RECT 1912.020 1017.370 1915.020 1017.380 ;
        RECT 2092.020 1017.370 2095.020 1017.380 ;
        RECT 2272.020 1017.370 2275.020 1017.380 ;
        RECT 2452.020 1017.370 2455.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.700 1017.370 2943.700 1017.380 ;
        RECT -24.080 840.380 -21.080 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1552.020 840.380 1555.020 840.390 ;
        RECT 1732.020 840.380 1735.020 840.390 ;
        RECT 1912.020 840.380 1915.020 840.390 ;
        RECT 2092.020 840.380 2095.020 840.390 ;
        RECT 2272.020 840.380 2275.020 840.390 ;
        RECT 2452.020 840.380 2455.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.700 840.380 2943.700 840.390 ;
        RECT -24.080 837.380 2943.700 840.380 ;
        RECT -24.080 837.370 -21.080 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1552.020 837.370 1555.020 837.380 ;
        RECT 1732.020 837.370 1735.020 837.380 ;
        RECT 1912.020 837.370 1915.020 837.380 ;
        RECT 2092.020 837.370 2095.020 837.380 ;
        RECT 2272.020 837.370 2275.020 837.380 ;
        RECT 2452.020 837.370 2455.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.700 837.370 2943.700 837.380 ;
        RECT -24.080 660.380 -21.080 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1552.020 660.380 1555.020 660.390 ;
        RECT 1732.020 660.380 1735.020 660.390 ;
        RECT 1912.020 660.380 1915.020 660.390 ;
        RECT 2092.020 660.380 2095.020 660.390 ;
        RECT 2272.020 660.380 2275.020 660.390 ;
        RECT 2452.020 660.380 2455.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.700 660.380 2943.700 660.390 ;
        RECT -24.080 657.380 2943.700 660.380 ;
        RECT -24.080 657.370 -21.080 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1552.020 657.370 1555.020 657.380 ;
        RECT 1732.020 657.370 1735.020 657.380 ;
        RECT 1912.020 657.370 1915.020 657.380 ;
        RECT 2092.020 657.370 2095.020 657.380 ;
        RECT 2272.020 657.370 2275.020 657.380 ;
        RECT 2452.020 657.370 2455.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.700 657.370 2943.700 657.380 ;
        RECT -24.080 480.380 -21.080 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.700 480.380 2943.700 480.390 ;
        RECT -24.080 477.380 2943.700 480.380 ;
        RECT -24.080 477.370 -21.080 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.700 477.370 2943.700 477.380 ;
        RECT -24.080 300.380 -21.080 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.700 300.380 2943.700 300.390 ;
        RECT -24.080 297.380 2943.700 300.380 ;
        RECT -24.080 297.370 -21.080 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.700 297.370 2943.700 297.380 ;
        RECT -24.080 120.380 -21.080 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.700 120.380 2943.700 120.390 ;
        RECT -24.080 117.380 2943.700 120.380 ;
        RECT -24.080 117.370 -21.080 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.700 117.370 2943.700 117.380 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 112.020 -15.720 115.020 -15.710 ;
        RECT 292.020 -15.720 295.020 -15.710 ;
        RECT 472.020 -15.720 475.020 -15.710 ;
        RECT 652.020 -15.720 655.020 -15.710 ;
        RECT 832.020 -15.720 835.020 -15.710 ;
        RECT 1012.020 -15.720 1015.020 -15.710 ;
        RECT 1192.020 -15.720 1195.020 -15.710 ;
        RECT 1372.020 -15.720 1375.020 -15.710 ;
        RECT 1552.020 -15.720 1555.020 -15.710 ;
        RECT 1732.020 -15.720 1735.020 -15.710 ;
        RECT 1912.020 -15.720 1915.020 -15.710 ;
        RECT 2092.020 -15.720 2095.020 -15.710 ;
        RECT 2272.020 -15.720 2275.020 -15.710 ;
        RECT 2452.020 -15.720 2455.020 -15.710 ;
        RECT 2632.020 -15.720 2635.020 -15.710 ;
        RECT 2812.020 -15.720 2815.020 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 112.020 -18.730 115.020 -18.720 ;
        RECT 292.020 -18.730 295.020 -18.720 ;
        RECT 472.020 -18.730 475.020 -18.720 ;
        RECT 652.020 -18.730 655.020 -18.720 ;
        RECT 832.020 -18.730 835.020 -18.720 ;
        RECT 1012.020 -18.730 1015.020 -18.720 ;
        RECT 1192.020 -18.730 1195.020 -18.720 ;
        RECT 1372.020 -18.730 1375.020 -18.720 ;
        RECT 1552.020 -18.730 1555.020 -18.720 ;
        RECT 1732.020 -18.730 1735.020 -18.720 ;
        RECT 1912.020 -18.730 1915.020 -18.720 ;
        RECT 2092.020 -18.730 2095.020 -18.720 ;
        RECT 2272.020 -18.730 2275.020 -18.720 ;
        RECT 2452.020 -18.730 2455.020 -18.720 ;
        RECT 2632.020 -18.730 2635.020 -18.720 ;
        RECT 2812.020 -18.730 2815.020 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT 40.020 -28.120 43.020 3547.800 ;
        RECT 220.020 -28.120 223.020 3547.800 ;
        RECT 400.020 -28.120 403.020 3547.800 ;
        RECT 580.020 -28.120 583.020 3547.800 ;
        RECT 760.020 -28.120 763.020 3547.800 ;
        RECT 940.020 -28.120 943.020 3547.800 ;
        RECT 1120.020 -28.120 1123.020 3547.800 ;
        RECT 1300.020 -28.120 1303.020 3547.800 ;
        RECT 1480.020 -28.120 1483.020 3547.800 ;
        RECT 1660.020 -28.120 1663.020 3547.800 ;
        RECT 1840.020 -28.120 1843.020 3547.800 ;
        RECT 2020.020 -28.120 2023.020 3547.800 ;
        RECT 2200.020 -28.120 2203.020 3547.800 ;
        RECT 2380.020 -28.120 2383.020 3547.800 ;
        RECT 2560.020 -28.120 2563.020 3547.800 ;
        RECT 2740.020 -28.120 2743.020 3547.800 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
      LAYER via4 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT -27.870 3467.090 -26.690 3468.270 ;
        RECT -27.870 3465.490 -26.690 3466.670 ;
        RECT -27.870 3287.090 -26.690 3288.270 ;
        RECT -27.870 3285.490 -26.690 3286.670 ;
        RECT -27.870 3107.090 -26.690 3108.270 ;
        RECT -27.870 3105.490 -26.690 3106.670 ;
        RECT -27.870 2927.090 -26.690 2928.270 ;
        RECT -27.870 2925.490 -26.690 2926.670 ;
        RECT -27.870 2747.090 -26.690 2748.270 ;
        RECT -27.870 2745.490 -26.690 2746.670 ;
        RECT -27.870 2567.090 -26.690 2568.270 ;
        RECT -27.870 2565.490 -26.690 2566.670 ;
        RECT -27.870 2387.090 -26.690 2388.270 ;
        RECT -27.870 2385.490 -26.690 2386.670 ;
        RECT -27.870 2207.090 -26.690 2208.270 ;
        RECT -27.870 2205.490 -26.690 2206.670 ;
        RECT -27.870 2027.090 -26.690 2028.270 ;
        RECT -27.870 2025.490 -26.690 2026.670 ;
        RECT -27.870 1847.090 -26.690 1848.270 ;
        RECT -27.870 1845.490 -26.690 1846.670 ;
        RECT -27.870 1667.090 -26.690 1668.270 ;
        RECT -27.870 1665.490 -26.690 1666.670 ;
        RECT -27.870 1487.090 -26.690 1488.270 ;
        RECT -27.870 1485.490 -26.690 1486.670 ;
        RECT -27.870 1307.090 -26.690 1308.270 ;
        RECT -27.870 1305.490 -26.690 1306.670 ;
        RECT -27.870 1127.090 -26.690 1128.270 ;
        RECT -27.870 1125.490 -26.690 1126.670 ;
        RECT -27.870 947.090 -26.690 948.270 ;
        RECT -27.870 945.490 -26.690 946.670 ;
        RECT -27.870 767.090 -26.690 768.270 ;
        RECT -27.870 765.490 -26.690 766.670 ;
        RECT -27.870 587.090 -26.690 588.270 ;
        RECT -27.870 585.490 -26.690 586.670 ;
        RECT -27.870 407.090 -26.690 408.270 ;
        RECT -27.870 405.490 -26.690 406.670 ;
        RECT -27.870 227.090 -26.690 228.270 ;
        RECT -27.870 225.490 -26.690 226.670 ;
        RECT -27.870 47.090 -26.690 48.270 ;
        RECT -27.870 45.490 -26.690 46.670 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 40.930 3541.810 42.110 3542.990 ;
        RECT 40.930 3540.210 42.110 3541.390 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.710 42.110 -20.530 ;
        RECT 40.930 -23.310 42.110 -22.130 ;
        RECT 220.930 3541.810 222.110 3542.990 ;
        RECT 220.930 3540.210 222.110 3541.390 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.710 222.110 -20.530 ;
        RECT 220.930 -23.310 222.110 -22.130 ;
        RECT 400.930 3541.810 402.110 3542.990 ;
        RECT 400.930 3540.210 402.110 3541.390 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 400.930 3107.090 402.110 3108.270 ;
        RECT 400.930 3105.490 402.110 3106.670 ;
        RECT 400.930 2927.090 402.110 2928.270 ;
        RECT 400.930 2925.490 402.110 2926.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 400.930 2567.090 402.110 2568.270 ;
        RECT 400.930 2565.490 402.110 2566.670 ;
        RECT 400.930 2387.090 402.110 2388.270 ;
        RECT 400.930 2385.490 402.110 2386.670 ;
        RECT 400.930 2207.090 402.110 2208.270 ;
        RECT 400.930 2205.490 402.110 2206.670 ;
        RECT 400.930 2027.090 402.110 2028.270 ;
        RECT 400.930 2025.490 402.110 2026.670 ;
        RECT 400.930 1847.090 402.110 1848.270 ;
        RECT 400.930 1845.490 402.110 1846.670 ;
        RECT 400.930 1667.090 402.110 1668.270 ;
        RECT 400.930 1665.490 402.110 1666.670 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.710 402.110 -20.530 ;
        RECT 400.930 -23.310 402.110 -22.130 ;
        RECT 580.930 3541.810 582.110 3542.990 ;
        RECT 580.930 3540.210 582.110 3541.390 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 580.930 3107.090 582.110 3108.270 ;
        RECT 580.930 3105.490 582.110 3106.670 ;
        RECT 580.930 2927.090 582.110 2928.270 ;
        RECT 580.930 2925.490 582.110 2926.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 580.930 2567.090 582.110 2568.270 ;
        RECT 580.930 2565.490 582.110 2566.670 ;
        RECT 580.930 2387.090 582.110 2388.270 ;
        RECT 580.930 2385.490 582.110 2386.670 ;
        RECT 580.930 2207.090 582.110 2208.270 ;
        RECT 580.930 2205.490 582.110 2206.670 ;
        RECT 580.930 2027.090 582.110 2028.270 ;
        RECT 580.930 2025.490 582.110 2026.670 ;
        RECT 580.930 1847.090 582.110 1848.270 ;
        RECT 580.930 1845.490 582.110 1846.670 ;
        RECT 580.930 1667.090 582.110 1668.270 ;
        RECT 580.930 1665.490 582.110 1666.670 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.710 582.110 -20.530 ;
        RECT 580.930 -23.310 582.110 -22.130 ;
        RECT 760.930 3541.810 762.110 3542.990 ;
        RECT 760.930 3540.210 762.110 3541.390 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 760.930 2567.090 762.110 2568.270 ;
        RECT 760.930 2565.490 762.110 2566.670 ;
        RECT 760.930 2387.090 762.110 2388.270 ;
        RECT 760.930 2385.490 762.110 2386.670 ;
        RECT 760.930 2207.090 762.110 2208.270 ;
        RECT 760.930 2205.490 762.110 2206.670 ;
        RECT 760.930 2027.090 762.110 2028.270 ;
        RECT 760.930 2025.490 762.110 2026.670 ;
        RECT 760.930 1847.090 762.110 1848.270 ;
        RECT 760.930 1845.490 762.110 1846.670 ;
        RECT 760.930 1667.090 762.110 1668.270 ;
        RECT 760.930 1665.490 762.110 1666.670 ;
        RECT 760.930 1487.090 762.110 1488.270 ;
        RECT 760.930 1485.490 762.110 1486.670 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 760.930 947.090 762.110 948.270 ;
        RECT 760.930 945.490 762.110 946.670 ;
        RECT 760.930 767.090 762.110 768.270 ;
        RECT 760.930 765.490 762.110 766.670 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.710 762.110 -20.530 ;
        RECT 760.930 -23.310 762.110 -22.130 ;
        RECT 940.930 3541.810 942.110 3542.990 ;
        RECT 940.930 3540.210 942.110 3541.390 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 940.930 2927.090 942.110 2928.270 ;
        RECT 940.930 2925.490 942.110 2926.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 940.930 2567.090 942.110 2568.270 ;
        RECT 940.930 2565.490 942.110 2566.670 ;
        RECT 940.930 2387.090 942.110 2388.270 ;
        RECT 940.930 2385.490 942.110 2386.670 ;
        RECT 940.930 2207.090 942.110 2208.270 ;
        RECT 940.930 2205.490 942.110 2206.670 ;
        RECT 940.930 2027.090 942.110 2028.270 ;
        RECT 940.930 2025.490 942.110 2026.670 ;
        RECT 940.930 1847.090 942.110 1848.270 ;
        RECT 940.930 1845.490 942.110 1846.670 ;
        RECT 940.930 1667.090 942.110 1668.270 ;
        RECT 940.930 1665.490 942.110 1666.670 ;
        RECT 940.930 1487.090 942.110 1488.270 ;
        RECT 940.930 1485.490 942.110 1486.670 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 940.930 947.090 942.110 948.270 ;
        RECT 940.930 945.490 942.110 946.670 ;
        RECT 940.930 767.090 942.110 768.270 ;
        RECT 940.930 765.490 942.110 766.670 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.710 942.110 -20.530 ;
        RECT 940.930 -23.310 942.110 -22.130 ;
        RECT 1120.930 3541.810 1122.110 3542.990 ;
        RECT 1120.930 3540.210 1122.110 3541.390 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1120.930 3107.090 1122.110 3108.270 ;
        RECT 1120.930 3105.490 1122.110 3106.670 ;
        RECT 1120.930 2927.090 1122.110 2928.270 ;
        RECT 1120.930 2925.490 1122.110 2926.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1120.930 2567.090 1122.110 2568.270 ;
        RECT 1120.930 2565.490 1122.110 2566.670 ;
        RECT 1120.930 2387.090 1122.110 2388.270 ;
        RECT 1120.930 2385.490 1122.110 2386.670 ;
        RECT 1120.930 2207.090 1122.110 2208.270 ;
        RECT 1120.930 2205.490 1122.110 2206.670 ;
        RECT 1120.930 2027.090 1122.110 2028.270 ;
        RECT 1120.930 2025.490 1122.110 2026.670 ;
        RECT 1120.930 1847.090 1122.110 1848.270 ;
        RECT 1120.930 1845.490 1122.110 1846.670 ;
        RECT 1120.930 1667.090 1122.110 1668.270 ;
        RECT 1120.930 1665.490 1122.110 1666.670 ;
        RECT 1120.930 1487.090 1122.110 1488.270 ;
        RECT 1120.930 1485.490 1122.110 1486.670 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1120.930 947.090 1122.110 948.270 ;
        RECT 1120.930 945.490 1122.110 946.670 ;
        RECT 1120.930 767.090 1122.110 768.270 ;
        RECT 1120.930 765.490 1122.110 766.670 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.710 1122.110 -20.530 ;
        RECT 1120.930 -23.310 1122.110 -22.130 ;
        RECT 1300.930 3541.810 1302.110 3542.990 ;
        RECT 1300.930 3540.210 1302.110 3541.390 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1300.930 3107.090 1302.110 3108.270 ;
        RECT 1300.930 3105.490 1302.110 3106.670 ;
        RECT 1300.930 2927.090 1302.110 2928.270 ;
        RECT 1300.930 2925.490 1302.110 2926.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1300.930 2567.090 1302.110 2568.270 ;
        RECT 1300.930 2565.490 1302.110 2566.670 ;
        RECT 1300.930 2387.090 1302.110 2388.270 ;
        RECT 1300.930 2385.490 1302.110 2386.670 ;
        RECT 1300.930 2207.090 1302.110 2208.270 ;
        RECT 1300.930 2205.490 1302.110 2206.670 ;
        RECT 1300.930 2027.090 1302.110 2028.270 ;
        RECT 1300.930 2025.490 1302.110 2026.670 ;
        RECT 1300.930 1847.090 1302.110 1848.270 ;
        RECT 1300.930 1845.490 1302.110 1846.670 ;
        RECT 1300.930 1667.090 1302.110 1668.270 ;
        RECT 1300.930 1665.490 1302.110 1666.670 ;
        RECT 1300.930 1487.090 1302.110 1488.270 ;
        RECT 1300.930 1485.490 1302.110 1486.670 ;
        RECT 1300.930 1307.090 1302.110 1308.270 ;
        RECT 1300.930 1305.490 1302.110 1306.670 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1300.930 947.090 1302.110 948.270 ;
        RECT 1300.930 945.490 1302.110 946.670 ;
        RECT 1300.930 767.090 1302.110 768.270 ;
        RECT 1300.930 765.490 1302.110 766.670 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.710 1302.110 -20.530 ;
        RECT 1300.930 -23.310 1302.110 -22.130 ;
        RECT 1480.930 3541.810 1482.110 3542.990 ;
        RECT 1480.930 3540.210 1482.110 3541.390 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 1480.930 2387.090 1482.110 2388.270 ;
        RECT 1480.930 2385.490 1482.110 2386.670 ;
        RECT 1480.930 2207.090 1482.110 2208.270 ;
        RECT 1480.930 2205.490 1482.110 2206.670 ;
        RECT 1480.930 2027.090 1482.110 2028.270 ;
        RECT 1480.930 2025.490 1482.110 2026.670 ;
        RECT 1480.930 1847.090 1482.110 1848.270 ;
        RECT 1480.930 1845.490 1482.110 1846.670 ;
        RECT 1480.930 1667.090 1482.110 1668.270 ;
        RECT 1480.930 1665.490 1482.110 1666.670 ;
        RECT 1480.930 1487.090 1482.110 1488.270 ;
        RECT 1480.930 1485.490 1482.110 1486.670 ;
        RECT 1480.930 1307.090 1482.110 1308.270 ;
        RECT 1480.930 1305.490 1482.110 1306.670 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1480.930 947.090 1482.110 948.270 ;
        RECT 1480.930 945.490 1482.110 946.670 ;
        RECT 1480.930 767.090 1482.110 768.270 ;
        RECT 1480.930 765.490 1482.110 766.670 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.710 1482.110 -20.530 ;
        RECT 1480.930 -23.310 1482.110 -22.130 ;
        RECT 1660.930 3541.810 1662.110 3542.990 ;
        RECT 1660.930 3540.210 1662.110 3541.390 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1660.930 2927.090 1662.110 2928.270 ;
        RECT 1660.930 2925.490 1662.110 2926.670 ;
        RECT 1660.930 2747.090 1662.110 2748.270 ;
        RECT 1660.930 2745.490 1662.110 2746.670 ;
        RECT 1660.930 2567.090 1662.110 2568.270 ;
        RECT 1660.930 2565.490 1662.110 2566.670 ;
        RECT 1660.930 2387.090 1662.110 2388.270 ;
        RECT 1660.930 2385.490 1662.110 2386.670 ;
        RECT 1660.930 2207.090 1662.110 2208.270 ;
        RECT 1660.930 2205.490 1662.110 2206.670 ;
        RECT 1660.930 2027.090 1662.110 2028.270 ;
        RECT 1660.930 2025.490 1662.110 2026.670 ;
        RECT 1660.930 1847.090 1662.110 1848.270 ;
        RECT 1660.930 1845.490 1662.110 1846.670 ;
        RECT 1660.930 1667.090 1662.110 1668.270 ;
        RECT 1660.930 1665.490 1662.110 1666.670 ;
        RECT 1660.930 1487.090 1662.110 1488.270 ;
        RECT 1660.930 1485.490 1662.110 1486.670 ;
        RECT 1660.930 1307.090 1662.110 1308.270 ;
        RECT 1660.930 1305.490 1662.110 1306.670 ;
        RECT 1660.930 1127.090 1662.110 1128.270 ;
        RECT 1660.930 1125.490 1662.110 1126.670 ;
        RECT 1660.930 947.090 1662.110 948.270 ;
        RECT 1660.930 945.490 1662.110 946.670 ;
        RECT 1660.930 767.090 1662.110 768.270 ;
        RECT 1660.930 765.490 1662.110 766.670 ;
        RECT 1660.930 587.090 1662.110 588.270 ;
        RECT 1660.930 585.490 1662.110 586.670 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.710 1662.110 -20.530 ;
        RECT 1660.930 -23.310 1662.110 -22.130 ;
        RECT 1840.930 3541.810 1842.110 3542.990 ;
        RECT 1840.930 3540.210 1842.110 3541.390 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 1840.930 2927.090 1842.110 2928.270 ;
        RECT 1840.930 2925.490 1842.110 2926.670 ;
        RECT 1840.930 2747.090 1842.110 2748.270 ;
        RECT 1840.930 2745.490 1842.110 2746.670 ;
        RECT 1840.930 2567.090 1842.110 2568.270 ;
        RECT 1840.930 2565.490 1842.110 2566.670 ;
        RECT 1840.930 2387.090 1842.110 2388.270 ;
        RECT 1840.930 2385.490 1842.110 2386.670 ;
        RECT 1840.930 2207.090 1842.110 2208.270 ;
        RECT 1840.930 2205.490 1842.110 2206.670 ;
        RECT 1840.930 2027.090 1842.110 2028.270 ;
        RECT 1840.930 2025.490 1842.110 2026.670 ;
        RECT 1840.930 1847.090 1842.110 1848.270 ;
        RECT 1840.930 1845.490 1842.110 1846.670 ;
        RECT 1840.930 1667.090 1842.110 1668.270 ;
        RECT 1840.930 1665.490 1842.110 1666.670 ;
        RECT 1840.930 1487.090 1842.110 1488.270 ;
        RECT 1840.930 1485.490 1842.110 1486.670 ;
        RECT 1840.930 1307.090 1842.110 1308.270 ;
        RECT 1840.930 1305.490 1842.110 1306.670 ;
        RECT 1840.930 1127.090 1842.110 1128.270 ;
        RECT 1840.930 1125.490 1842.110 1126.670 ;
        RECT 1840.930 947.090 1842.110 948.270 ;
        RECT 1840.930 945.490 1842.110 946.670 ;
        RECT 1840.930 767.090 1842.110 768.270 ;
        RECT 1840.930 765.490 1842.110 766.670 ;
        RECT 1840.930 587.090 1842.110 588.270 ;
        RECT 1840.930 585.490 1842.110 586.670 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.710 1842.110 -20.530 ;
        RECT 1840.930 -23.310 1842.110 -22.130 ;
        RECT 2020.930 3541.810 2022.110 3542.990 ;
        RECT 2020.930 3540.210 2022.110 3541.390 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 2020.930 2387.090 2022.110 2388.270 ;
        RECT 2020.930 2385.490 2022.110 2386.670 ;
        RECT 2020.930 2207.090 2022.110 2208.270 ;
        RECT 2020.930 2205.490 2022.110 2206.670 ;
        RECT 2020.930 2027.090 2022.110 2028.270 ;
        RECT 2020.930 2025.490 2022.110 2026.670 ;
        RECT 2020.930 1847.090 2022.110 1848.270 ;
        RECT 2020.930 1845.490 2022.110 1846.670 ;
        RECT 2020.930 1667.090 2022.110 1668.270 ;
        RECT 2020.930 1665.490 2022.110 1666.670 ;
        RECT 2020.930 1487.090 2022.110 1488.270 ;
        RECT 2020.930 1485.490 2022.110 1486.670 ;
        RECT 2020.930 1307.090 2022.110 1308.270 ;
        RECT 2020.930 1305.490 2022.110 1306.670 ;
        RECT 2020.930 1127.090 2022.110 1128.270 ;
        RECT 2020.930 1125.490 2022.110 1126.670 ;
        RECT 2020.930 947.090 2022.110 948.270 ;
        RECT 2020.930 945.490 2022.110 946.670 ;
        RECT 2020.930 767.090 2022.110 768.270 ;
        RECT 2020.930 765.490 2022.110 766.670 ;
        RECT 2020.930 587.090 2022.110 588.270 ;
        RECT 2020.930 585.490 2022.110 586.670 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.710 2022.110 -20.530 ;
        RECT 2020.930 -23.310 2022.110 -22.130 ;
        RECT 2200.930 3541.810 2202.110 3542.990 ;
        RECT 2200.930 3540.210 2202.110 3541.390 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2200.930 2927.090 2202.110 2928.270 ;
        RECT 2200.930 2925.490 2202.110 2926.670 ;
        RECT 2200.930 2747.090 2202.110 2748.270 ;
        RECT 2200.930 2745.490 2202.110 2746.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2200.930 2387.090 2202.110 2388.270 ;
        RECT 2200.930 2385.490 2202.110 2386.670 ;
        RECT 2200.930 2207.090 2202.110 2208.270 ;
        RECT 2200.930 2205.490 2202.110 2206.670 ;
        RECT 2200.930 2027.090 2202.110 2028.270 ;
        RECT 2200.930 2025.490 2202.110 2026.670 ;
        RECT 2200.930 1847.090 2202.110 1848.270 ;
        RECT 2200.930 1845.490 2202.110 1846.670 ;
        RECT 2200.930 1667.090 2202.110 1668.270 ;
        RECT 2200.930 1665.490 2202.110 1666.670 ;
        RECT 2200.930 1487.090 2202.110 1488.270 ;
        RECT 2200.930 1485.490 2202.110 1486.670 ;
        RECT 2200.930 1307.090 2202.110 1308.270 ;
        RECT 2200.930 1305.490 2202.110 1306.670 ;
        RECT 2200.930 1127.090 2202.110 1128.270 ;
        RECT 2200.930 1125.490 2202.110 1126.670 ;
        RECT 2200.930 947.090 2202.110 948.270 ;
        RECT 2200.930 945.490 2202.110 946.670 ;
        RECT 2200.930 767.090 2202.110 768.270 ;
        RECT 2200.930 765.490 2202.110 766.670 ;
        RECT 2200.930 587.090 2202.110 588.270 ;
        RECT 2200.930 585.490 2202.110 586.670 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.710 2202.110 -20.530 ;
        RECT 2200.930 -23.310 2202.110 -22.130 ;
        RECT 2380.930 3541.810 2382.110 3542.990 ;
        RECT 2380.930 3540.210 2382.110 3541.390 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2380.930 2927.090 2382.110 2928.270 ;
        RECT 2380.930 2925.490 2382.110 2926.670 ;
        RECT 2380.930 2747.090 2382.110 2748.270 ;
        RECT 2380.930 2745.490 2382.110 2746.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2380.930 2387.090 2382.110 2388.270 ;
        RECT 2380.930 2385.490 2382.110 2386.670 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2380.930 2027.090 2382.110 2028.270 ;
        RECT 2380.930 2025.490 2382.110 2026.670 ;
        RECT 2380.930 1847.090 2382.110 1848.270 ;
        RECT 2380.930 1845.490 2382.110 1846.670 ;
        RECT 2380.930 1667.090 2382.110 1668.270 ;
        RECT 2380.930 1665.490 2382.110 1666.670 ;
        RECT 2380.930 1487.090 2382.110 1488.270 ;
        RECT 2380.930 1485.490 2382.110 1486.670 ;
        RECT 2380.930 1307.090 2382.110 1308.270 ;
        RECT 2380.930 1305.490 2382.110 1306.670 ;
        RECT 2380.930 1127.090 2382.110 1128.270 ;
        RECT 2380.930 1125.490 2382.110 1126.670 ;
        RECT 2380.930 947.090 2382.110 948.270 ;
        RECT 2380.930 945.490 2382.110 946.670 ;
        RECT 2380.930 767.090 2382.110 768.270 ;
        RECT 2380.930 765.490 2382.110 766.670 ;
        RECT 2380.930 587.090 2382.110 588.270 ;
        RECT 2380.930 585.490 2382.110 586.670 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.710 2382.110 -20.530 ;
        RECT 2380.930 -23.310 2382.110 -22.130 ;
        RECT 2560.930 3541.810 2562.110 3542.990 ;
        RECT 2560.930 3540.210 2562.110 3541.390 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.710 2562.110 -20.530 ;
        RECT 2560.930 -23.310 2562.110 -22.130 ;
        RECT 2740.930 3541.810 2742.110 3542.990 ;
        RECT 2740.930 3540.210 2742.110 3541.390 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.710 2742.110 -20.530 ;
        RECT 2740.930 -23.310 2742.110 -22.130 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT 2946.310 3467.090 2947.490 3468.270 ;
        RECT 2946.310 3465.490 2947.490 3466.670 ;
        RECT 2946.310 3287.090 2947.490 3288.270 ;
        RECT 2946.310 3285.490 2947.490 3286.670 ;
        RECT 2946.310 3107.090 2947.490 3108.270 ;
        RECT 2946.310 3105.490 2947.490 3106.670 ;
        RECT 2946.310 2927.090 2947.490 2928.270 ;
        RECT 2946.310 2925.490 2947.490 2926.670 ;
        RECT 2946.310 2747.090 2947.490 2748.270 ;
        RECT 2946.310 2745.490 2947.490 2746.670 ;
        RECT 2946.310 2567.090 2947.490 2568.270 ;
        RECT 2946.310 2565.490 2947.490 2566.670 ;
        RECT 2946.310 2387.090 2947.490 2388.270 ;
        RECT 2946.310 2385.490 2947.490 2386.670 ;
        RECT 2946.310 2207.090 2947.490 2208.270 ;
        RECT 2946.310 2205.490 2947.490 2206.670 ;
        RECT 2946.310 2027.090 2947.490 2028.270 ;
        RECT 2946.310 2025.490 2947.490 2026.670 ;
        RECT 2946.310 1847.090 2947.490 1848.270 ;
        RECT 2946.310 1845.490 2947.490 1846.670 ;
        RECT 2946.310 1667.090 2947.490 1668.270 ;
        RECT 2946.310 1665.490 2947.490 1666.670 ;
        RECT 2946.310 1487.090 2947.490 1488.270 ;
        RECT 2946.310 1485.490 2947.490 1486.670 ;
        RECT 2946.310 1307.090 2947.490 1308.270 ;
        RECT 2946.310 1305.490 2947.490 1306.670 ;
        RECT 2946.310 1127.090 2947.490 1128.270 ;
        RECT 2946.310 1125.490 2947.490 1126.670 ;
        RECT 2946.310 947.090 2947.490 948.270 ;
        RECT 2946.310 945.490 2947.490 946.670 ;
        RECT 2946.310 767.090 2947.490 768.270 ;
        RECT 2946.310 765.490 2947.490 766.670 ;
        RECT 2946.310 587.090 2947.490 588.270 ;
        RECT 2946.310 585.490 2947.490 586.670 ;
        RECT 2946.310 407.090 2947.490 408.270 ;
        RECT 2946.310 405.490 2947.490 406.670 ;
        RECT 2946.310 227.090 2947.490 228.270 ;
        RECT 2946.310 225.490 2947.490 226.670 ;
        RECT 2946.310 47.090 2947.490 48.270 ;
        RECT 2946.310 45.490 2947.490 46.670 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
      LAYER met5 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 40.020 3543.100 43.020 3543.110 ;
        RECT 220.020 3543.100 223.020 3543.110 ;
        RECT 400.020 3543.100 403.020 3543.110 ;
        RECT 580.020 3543.100 583.020 3543.110 ;
        RECT 760.020 3543.100 763.020 3543.110 ;
        RECT 940.020 3543.100 943.020 3543.110 ;
        RECT 1120.020 3543.100 1123.020 3543.110 ;
        RECT 1300.020 3543.100 1303.020 3543.110 ;
        RECT 1480.020 3543.100 1483.020 3543.110 ;
        RECT 1660.020 3543.100 1663.020 3543.110 ;
        RECT 1840.020 3543.100 1843.020 3543.110 ;
        RECT 2020.020 3543.100 2023.020 3543.110 ;
        RECT 2200.020 3543.100 2203.020 3543.110 ;
        RECT 2380.020 3543.100 2383.020 3543.110 ;
        RECT 2560.020 3543.100 2563.020 3543.110 ;
        RECT 2740.020 3543.100 2743.020 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 40.020 3540.090 43.020 3540.100 ;
        RECT 220.020 3540.090 223.020 3540.100 ;
        RECT 400.020 3540.090 403.020 3540.100 ;
        RECT 580.020 3540.090 583.020 3540.100 ;
        RECT 760.020 3540.090 763.020 3540.100 ;
        RECT 940.020 3540.090 943.020 3540.100 ;
        RECT 1120.020 3540.090 1123.020 3540.100 ;
        RECT 1300.020 3540.090 1303.020 3540.100 ;
        RECT 1480.020 3540.090 1483.020 3540.100 ;
        RECT 1660.020 3540.090 1663.020 3540.100 ;
        RECT 1840.020 3540.090 1843.020 3540.100 ;
        RECT 2020.020 3540.090 2023.020 3540.100 ;
        RECT 2200.020 3540.090 2203.020 3540.100 ;
        RECT 2380.020 3540.090 2383.020 3540.100 ;
        RECT 2560.020 3540.090 2563.020 3540.100 ;
        RECT 2740.020 3540.090 2743.020 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -28.780 3468.380 -25.780 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.400 3468.380 2948.400 3468.390 ;
        RECT -33.480 3465.380 2953.100 3468.380 ;
        RECT -28.780 3465.370 -25.780 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.400 3465.370 2948.400 3465.380 ;
        RECT -28.780 3288.380 -25.780 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.400 3288.380 2948.400 3288.390 ;
        RECT -33.480 3285.380 2953.100 3288.380 ;
        RECT -28.780 3285.370 -25.780 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.400 3285.370 2948.400 3285.380 ;
        RECT -28.780 3108.380 -25.780 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 400.020 3108.380 403.020 3108.390 ;
        RECT 580.020 3108.380 583.020 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1120.020 3108.380 1123.020 3108.390 ;
        RECT 1300.020 3108.380 1303.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.400 3108.380 2948.400 3108.390 ;
        RECT -33.480 3105.380 2953.100 3108.380 ;
        RECT -28.780 3105.370 -25.780 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 400.020 3105.370 403.020 3105.380 ;
        RECT 580.020 3105.370 583.020 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1120.020 3105.370 1123.020 3105.380 ;
        RECT 1300.020 3105.370 1303.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.400 3105.370 2948.400 3105.380 ;
        RECT -28.780 2928.380 -25.780 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 400.020 2928.380 403.020 2928.390 ;
        RECT 580.020 2928.380 583.020 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 940.020 2928.380 943.020 2928.390 ;
        RECT 1120.020 2928.380 1123.020 2928.390 ;
        RECT 1300.020 2928.380 1303.020 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1660.020 2928.380 1663.020 2928.390 ;
        RECT 1840.020 2928.380 1843.020 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2200.020 2928.380 2203.020 2928.390 ;
        RECT 2380.020 2928.380 2383.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.400 2928.380 2948.400 2928.390 ;
        RECT -33.480 2925.380 2953.100 2928.380 ;
        RECT -28.780 2925.370 -25.780 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 400.020 2925.370 403.020 2925.380 ;
        RECT 580.020 2925.370 583.020 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 940.020 2925.370 943.020 2925.380 ;
        RECT 1120.020 2925.370 1123.020 2925.380 ;
        RECT 1300.020 2925.370 1303.020 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1660.020 2925.370 1663.020 2925.380 ;
        RECT 1840.020 2925.370 1843.020 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2200.020 2925.370 2203.020 2925.380 ;
        RECT 2380.020 2925.370 2383.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.400 2925.370 2948.400 2925.380 ;
        RECT -28.780 2748.380 -25.780 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 1660.020 2748.380 1663.020 2748.390 ;
        RECT 1840.020 2748.380 1843.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2200.020 2748.380 2203.020 2748.390 ;
        RECT 2380.020 2748.380 2383.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.400 2748.380 2948.400 2748.390 ;
        RECT -33.480 2745.380 2953.100 2748.380 ;
        RECT -28.780 2745.370 -25.780 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 1660.020 2745.370 1663.020 2745.380 ;
        RECT 1840.020 2745.370 1843.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2200.020 2745.370 2203.020 2745.380 ;
        RECT 2380.020 2745.370 2383.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.400 2745.370 2948.400 2745.380 ;
        RECT -28.780 2568.380 -25.780 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 400.020 2568.380 403.020 2568.390 ;
        RECT 580.020 2568.380 583.020 2568.390 ;
        RECT 760.020 2568.380 763.020 2568.390 ;
        RECT 940.020 2568.380 943.020 2568.390 ;
        RECT 1120.020 2568.380 1123.020 2568.390 ;
        RECT 1300.020 2568.380 1303.020 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 1660.020 2568.380 1663.020 2568.390 ;
        RECT 1840.020 2568.380 1843.020 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.400 2568.380 2948.400 2568.390 ;
        RECT -33.480 2565.380 2953.100 2568.380 ;
        RECT -28.780 2565.370 -25.780 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 400.020 2565.370 403.020 2565.380 ;
        RECT 580.020 2565.370 583.020 2565.380 ;
        RECT 760.020 2565.370 763.020 2565.380 ;
        RECT 940.020 2565.370 943.020 2565.380 ;
        RECT 1120.020 2565.370 1123.020 2565.380 ;
        RECT 1300.020 2565.370 1303.020 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 1660.020 2565.370 1663.020 2565.380 ;
        RECT 1840.020 2565.370 1843.020 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.400 2565.370 2948.400 2565.380 ;
        RECT -28.780 2388.380 -25.780 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 400.020 2388.380 403.020 2388.390 ;
        RECT 580.020 2388.380 583.020 2388.390 ;
        RECT 760.020 2388.380 763.020 2388.390 ;
        RECT 940.020 2388.380 943.020 2388.390 ;
        RECT 1120.020 2388.380 1123.020 2388.390 ;
        RECT 1300.020 2388.380 1303.020 2388.390 ;
        RECT 1480.020 2388.380 1483.020 2388.390 ;
        RECT 1660.020 2388.380 1663.020 2388.390 ;
        RECT 1840.020 2388.380 1843.020 2388.390 ;
        RECT 2020.020 2388.380 2023.020 2388.390 ;
        RECT 2200.020 2388.380 2203.020 2388.390 ;
        RECT 2380.020 2388.380 2383.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.400 2388.380 2948.400 2388.390 ;
        RECT -33.480 2385.380 2953.100 2388.380 ;
        RECT -28.780 2385.370 -25.780 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 400.020 2385.370 403.020 2385.380 ;
        RECT 580.020 2385.370 583.020 2385.380 ;
        RECT 760.020 2385.370 763.020 2385.380 ;
        RECT 940.020 2385.370 943.020 2385.380 ;
        RECT 1120.020 2385.370 1123.020 2385.380 ;
        RECT 1300.020 2385.370 1303.020 2385.380 ;
        RECT 1480.020 2385.370 1483.020 2385.380 ;
        RECT 1660.020 2385.370 1663.020 2385.380 ;
        RECT 1840.020 2385.370 1843.020 2385.380 ;
        RECT 2020.020 2385.370 2023.020 2385.380 ;
        RECT 2200.020 2385.370 2203.020 2385.380 ;
        RECT 2380.020 2385.370 2383.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.400 2385.370 2948.400 2385.380 ;
        RECT -28.780 2208.380 -25.780 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 400.020 2208.380 403.020 2208.390 ;
        RECT 580.020 2208.380 583.020 2208.390 ;
        RECT 760.020 2208.380 763.020 2208.390 ;
        RECT 940.020 2208.380 943.020 2208.390 ;
        RECT 1120.020 2208.380 1123.020 2208.390 ;
        RECT 1300.020 2208.380 1303.020 2208.390 ;
        RECT 1480.020 2208.380 1483.020 2208.390 ;
        RECT 1660.020 2208.380 1663.020 2208.390 ;
        RECT 1840.020 2208.380 1843.020 2208.390 ;
        RECT 2020.020 2208.380 2023.020 2208.390 ;
        RECT 2200.020 2208.380 2203.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.400 2208.380 2948.400 2208.390 ;
        RECT -33.480 2205.380 2953.100 2208.380 ;
        RECT -28.780 2205.370 -25.780 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 400.020 2205.370 403.020 2205.380 ;
        RECT 580.020 2205.370 583.020 2205.380 ;
        RECT 760.020 2205.370 763.020 2205.380 ;
        RECT 940.020 2205.370 943.020 2205.380 ;
        RECT 1120.020 2205.370 1123.020 2205.380 ;
        RECT 1300.020 2205.370 1303.020 2205.380 ;
        RECT 1480.020 2205.370 1483.020 2205.380 ;
        RECT 1660.020 2205.370 1663.020 2205.380 ;
        RECT 1840.020 2205.370 1843.020 2205.380 ;
        RECT 2020.020 2205.370 2023.020 2205.380 ;
        RECT 2200.020 2205.370 2203.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.400 2205.370 2948.400 2205.380 ;
        RECT -28.780 2028.380 -25.780 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 400.020 2028.380 403.020 2028.390 ;
        RECT 580.020 2028.380 583.020 2028.390 ;
        RECT 760.020 2028.380 763.020 2028.390 ;
        RECT 940.020 2028.380 943.020 2028.390 ;
        RECT 1120.020 2028.380 1123.020 2028.390 ;
        RECT 1300.020 2028.380 1303.020 2028.390 ;
        RECT 1480.020 2028.380 1483.020 2028.390 ;
        RECT 1660.020 2028.380 1663.020 2028.390 ;
        RECT 1840.020 2028.380 1843.020 2028.390 ;
        RECT 2020.020 2028.380 2023.020 2028.390 ;
        RECT 2200.020 2028.380 2203.020 2028.390 ;
        RECT 2380.020 2028.380 2383.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.400 2028.380 2948.400 2028.390 ;
        RECT -33.480 2025.380 2953.100 2028.380 ;
        RECT -28.780 2025.370 -25.780 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 400.020 2025.370 403.020 2025.380 ;
        RECT 580.020 2025.370 583.020 2025.380 ;
        RECT 760.020 2025.370 763.020 2025.380 ;
        RECT 940.020 2025.370 943.020 2025.380 ;
        RECT 1120.020 2025.370 1123.020 2025.380 ;
        RECT 1300.020 2025.370 1303.020 2025.380 ;
        RECT 1480.020 2025.370 1483.020 2025.380 ;
        RECT 1660.020 2025.370 1663.020 2025.380 ;
        RECT 1840.020 2025.370 1843.020 2025.380 ;
        RECT 2020.020 2025.370 2023.020 2025.380 ;
        RECT 2200.020 2025.370 2203.020 2025.380 ;
        RECT 2380.020 2025.370 2383.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.400 2025.370 2948.400 2025.380 ;
        RECT -28.780 1848.380 -25.780 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 400.020 1848.380 403.020 1848.390 ;
        RECT 580.020 1848.380 583.020 1848.390 ;
        RECT 760.020 1848.380 763.020 1848.390 ;
        RECT 940.020 1848.380 943.020 1848.390 ;
        RECT 1120.020 1848.380 1123.020 1848.390 ;
        RECT 1300.020 1848.380 1303.020 1848.390 ;
        RECT 1480.020 1848.380 1483.020 1848.390 ;
        RECT 1660.020 1848.380 1663.020 1848.390 ;
        RECT 1840.020 1848.380 1843.020 1848.390 ;
        RECT 2020.020 1848.380 2023.020 1848.390 ;
        RECT 2200.020 1848.380 2203.020 1848.390 ;
        RECT 2380.020 1848.380 2383.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.400 1848.380 2948.400 1848.390 ;
        RECT -33.480 1845.380 2953.100 1848.380 ;
        RECT -28.780 1845.370 -25.780 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 400.020 1845.370 403.020 1845.380 ;
        RECT 580.020 1845.370 583.020 1845.380 ;
        RECT 760.020 1845.370 763.020 1845.380 ;
        RECT 940.020 1845.370 943.020 1845.380 ;
        RECT 1120.020 1845.370 1123.020 1845.380 ;
        RECT 1300.020 1845.370 1303.020 1845.380 ;
        RECT 1480.020 1845.370 1483.020 1845.380 ;
        RECT 1660.020 1845.370 1663.020 1845.380 ;
        RECT 1840.020 1845.370 1843.020 1845.380 ;
        RECT 2020.020 1845.370 2023.020 1845.380 ;
        RECT 2200.020 1845.370 2203.020 1845.380 ;
        RECT 2380.020 1845.370 2383.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.400 1845.370 2948.400 1845.380 ;
        RECT -28.780 1668.380 -25.780 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 400.020 1668.380 403.020 1668.390 ;
        RECT 580.020 1668.380 583.020 1668.390 ;
        RECT 760.020 1668.380 763.020 1668.390 ;
        RECT 940.020 1668.380 943.020 1668.390 ;
        RECT 1120.020 1668.380 1123.020 1668.390 ;
        RECT 1300.020 1668.380 1303.020 1668.390 ;
        RECT 1480.020 1668.380 1483.020 1668.390 ;
        RECT 1660.020 1668.380 1663.020 1668.390 ;
        RECT 1840.020 1668.380 1843.020 1668.390 ;
        RECT 2020.020 1668.380 2023.020 1668.390 ;
        RECT 2200.020 1668.380 2203.020 1668.390 ;
        RECT 2380.020 1668.380 2383.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.400 1668.380 2948.400 1668.390 ;
        RECT -33.480 1665.380 2953.100 1668.380 ;
        RECT -28.780 1665.370 -25.780 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 400.020 1665.370 403.020 1665.380 ;
        RECT 580.020 1665.370 583.020 1665.380 ;
        RECT 760.020 1665.370 763.020 1665.380 ;
        RECT 940.020 1665.370 943.020 1665.380 ;
        RECT 1120.020 1665.370 1123.020 1665.380 ;
        RECT 1300.020 1665.370 1303.020 1665.380 ;
        RECT 1480.020 1665.370 1483.020 1665.380 ;
        RECT 1660.020 1665.370 1663.020 1665.380 ;
        RECT 1840.020 1665.370 1843.020 1665.380 ;
        RECT 2020.020 1665.370 2023.020 1665.380 ;
        RECT 2200.020 1665.370 2203.020 1665.380 ;
        RECT 2380.020 1665.370 2383.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.400 1665.370 2948.400 1665.380 ;
        RECT -28.780 1488.380 -25.780 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 760.020 1488.380 763.020 1488.390 ;
        RECT 940.020 1488.380 943.020 1488.390 ;
        RECT 1120.020 1488.380 1123.020 1488.390 ;
        RECT 1300.020 1488.380 1303.020 1488.390 ;
        RECT 1480.020 1488.380 1483.020 1488.390 ;
        RECT 1660.020 1488.380 1663.020 1488.390 ;
        RECT 1840.020 1488.380 1843.020 1488.390 ;
        RECT 2020.020 1488.380 2023.020 1488.390 ;
        RECT 2200.020 1488.380 2203.020 1488.390 ;
        RECT 2380.020 1488.380 2383.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.400 1488.380 2948.400 1488.390 ;
        RECT -33.480 1485.380 2953.100 1488.380 ;
        RECT -28.780 1485.370 -25.780 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 760.020 1485.370 763.020 1485.380 ;
        RECT 940.020 1485.370 943.020 1485.380 ;
        RECT 1120.020 1485.370 1123.020 1485.380 ;
        RECT 1300.020 1485.370 1303.020 1485.380 ;
        RECT 1480.020 1485.370 1483.020 1485.380 ;
        RECT 1660.020 1485.370 1663.020 1485.380 ;
        RECT 1840.020 1485.370 1843.020 1485.380 ;
        RECT 2020.020 1485.370 2023.020 1485.380 ;
        RECT 2200.020 1485.370 2203.020 1485.380 ;
        RECT 2380.020 1485.370 2383.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.400 1485.370 2948.400 1485.380 ;
        RECT -28.780 1308.380 -25.780 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 1300.020 1308.380 1303.020 1308.390 ;
        RECT 1480.020 1308.380 1483.020 1308.390 ;
        RECT 1660.020 1308.380 1663.020 1308.390 ;
        RECT 1840.020 1308.380 1843.020 1308.390 ;
        RECT 2020.020 1308.380 2023.020 1308.390 ;
        RECT 2200.020 1308.380 2203.020 1308.390 ;
        RECT 2380.020 1308.380 2383.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.400 1308.380 2948.400 1308.390 ;
        RECT -33.480 1305.380 2953.100 1308.380 ;
        RECT -28.780 1305.370 -25.780 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 1300.020 1305.370 1303.020 1305.380 ;
        RECT 1480.020 1305.370 1483.020 1305.380 ;
        RECT 1660.020 1305.370 1663.020 1305.380 ;
        RECT 1840.020 1305.370 1843.020 1305.380 ;
        RECT 2020.020 1305.370 2023.020 1305.380 ;
        RECT 2200.020 1305.370 2203.020 1305.380 ;
        RECT 2380.020 1305.370 2383.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.400 1305.370 2948.400 1305.380 ;
        RECT -28.780 1128.380 -25.780 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1660.020 1128.380 1663.020 1128.390 ;
        RECT 1840.020 1128.380 1843.020 1128.390 ;
        RECT 2020.020 1128.380 2023.020 1128.390 ;
        RECT 2200.020 1128.380 2203.020 1128.390 ;
        RECT 2380.020 1128.380 2383.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.400 1128.380 2948.400 1128.390 ;
        RECT -33.480 1125.380 2953.100 1128.380 ;
        RECT -28.780 1125.370 -25.780 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1660.020 1125.370 1663.020 1125.380 ;
        RECT 1840.020 1125.370 1843.020 1125.380 ;
        RECT 2020.020 1125.370 2023.020 1125.380 ;
        RECT 2200.020 1125.370 2203.020 1125.380 ;
        RECT 2380.020 1125.370 2383.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.400 1125.370 2948.400 1125.380 ;
        RECT -28.780 948.380 -25.780 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 760.020 948.380 763.020 948.390 ;
        RECT 940.020 948.380 943.020 948.390 ;
        RECT 1120.020 948.380 1123.020 948.390 ;
        RECT 1300.020 948.380 1303.020 948.390 ;
        RECT 1480.020 948.380 1483.020 948.390 ;
        RECT 1660.020 948.380 1663.020 948.390 ;
        RECT 1840.020 948.380 1843.020 948.390 ;
        RECT 2020.020 948.380 2023.020 948.390 ;
        RECT 2200.020 948.380 2203.020 948.390 ;
        RECT 2380.020 948.380 2383.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.400 948.380 2948.400 948.390 ;
        RECT -33.480 945.380 2953.100 948.380 ;
        RECT -28.780 945.370 -25.780 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 760.020 945.370 763.020 945.380 ;
        RECT 940.020 945.370 943.020 945.380 ;
        RECT 1120.020 945.370 1123.020 945.380 ;
        RECT 1300.020 945.370 1303.020 945.380 ;
        RECT 1480.020 945.370 1483.020 945.380 ;
        RECT 1660.020 945.370 1663.020 945.380 ;
        RECT 1840.020 945.370 1843.020 945.380 ;
        RECT 2020.020 945.370 2023.020 945.380 ;
        RECT 2200.020 945.370 2203.020 945.380 ;
        RECT 2380.020 945.370 2383.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.400 945.370 2948.400 945.380 ;
        RECT -28.780 768.380 -25.780 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 760.020 768.380 763.020 768.390 ;
        RECT 940.020 768.380 943.020 768.390 ;
        RECT 1120.020 768.380 1123.020 768.390 ;
        RECT 1300.020 768.380 1303.020 768.390 ;
        RECT 1480.020 768.380 1483.020 768.390 ;
        RECT 1660.020 768.380 1663.020 768.390 ;
        RECT 1840.020 768.380 1843.020 768.390 ;
        RECT 2020.020 768.380 2023.020 768.390 ;
        RECT 2200.020 768.380 2203.020 768.390 ;
        RECT 2380.020 768.380 2383.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.400 768.380 2948.400 768.390 ;
        RECT -33.480 765.380 2953.100 768.380 ;
        RECT -28.780 765.370 -25.780 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 760.020 765.370 763.020 765.380 ;
        RECT 940.020 765.370 943.020 765.380 ;
        RECT 1120.020 765.370 1123.020 765.380 ;
        RECT 1300.020 765.370 1303.020 765.380 ;
        RECT 1480.020 765.370 1483.020 765.380 ;
        RECT 1660.020 765.370 1663.020 765.380 ;
        RECT 1840.020 765.370 1843.020 765.380 ;
        RECT 2020.020 765.370 2023.020 765.380 ;
        RECT 2200.020 765.370 2203.020 765.380 ;
        RECT 2380.020 765.370 2383.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.400 765.370 2948.400 765.380 ;
        RECT -28.780 588.380 -25.780 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1660.020 588.380 1663.020 588.390 ;
        RECT 1840.020 588.380 1843.020 588.390 ;
        RECT 2020.020 588.380 2023.020 588.390 ;
        RECT 2200.020 588.380 2203.020 588.390 ;
        RECT 2380.020 588.380 2383.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.400 588.380 2948.400 588.390 ;
        RECT -33.480 585.380 2953.100 588.380 ;
        RECT -28.780 585.370 -25.780 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1660.020 585.370 1663.020 585.380 ;
        RECT 1840.020 585.370 1843.020 585.380 ;
        RECT 2020.020 585.370 2023.020 585.380 ;
        RECT 2200.020 585.370 2203.020 585.380 ;
        RECT 2380.020 585.370 2383.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.400 585.370 2948.400 585.380 ;
        RECT -28.780 408.380 -25.780 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.400 408.380 2948.400 408.390 ;
        RECT -33.480 405.380 2953.100 408.380 ;
        RECT -28.780 405.370 -25.780 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.400 405.370 2948.400 405.380 ;
        RECT -28.780 228.380 -25.780 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.400 228.380 2948.400 228.390 ;
        RECT -33.480 225.380 2953.100 228.380 ;
        RECT -28.780 225.370 -25.780 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.400 225.370 2948.400 225.380 ;
        RECT -28.780 48.380 -25.780 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.400 48.380 2948.400 48.390 ;
        RECT -33.480 45.380 2953.100 48.380 ;
        RECT -28.780 45.370 -25.780 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.400 45.370 2948.400 45.380 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 40.020 -20.420 43.020 -20.410 ;
        RECT 220.020 -20.420 223.020 -20.410 ;
        RECT 400.020 -20.420 403.020 -20.410 ;
        RECT 580.020 -20.420 583.020 -20.410 ;
        RECT 760.020 -20.420 763.020 -20.410 ;
        RECT 940.020 -20.420 943.020 -20.410 ;
        RECT 1120.020 -20.420 1123.020 -20.410 ;
        RECT 1300.020 -20.420 1303.020 -20.410 ;
        RECT 1480.020 -20.420 1483.020 -20.410 ;
        RECT 1660.020 -20.420 1663.020 -20.410 ;
        RECT 1840.020 -20.420 1843.020 -20.410 ;
        RECT 2020.020 -20.420 2023.020 -20.410 ;
        RECT 2200.020 -20.420 2203.020 -20.410 ;
        RECT 2380.020 -20.420 2383.020 -20.410 ;
        RECT 2560.020 -20.420 2563.020 -20.410 ;
        RECT 2740.020 -20.420 2743.020 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 40.020 -23.430 43.020 -23.420 ;
        RECT 220.020 -23.430 223.020 -23.420 ;
        RECT 400.020 -23.430 403.020 -23.420 ;
        RECT 580.020 -23.430 583.020 -23.420 ;
        RECT 760.020 -23.430 763.020 -23.420 ;
        RECT 940.020 -23.430 943.020 -23.420 ;
        RECT 1120.020 -23.430 1123.020 -23.420 ;
        RECT 1300.020 -23.430 1303.020 -23.420 ;
        RECT 1480.020 -23.430 1483.020 -23.420 ;
        RECT 1660.020 -23.430 1663.020 -23.420 ;
        RECT 1840.020 -23.430 1843.020 -23.420 ;
        RECT 2020.020 -23.430 2023.020 -23.420 ;
        RECT 2200.020 -23.430 2203.020 -23.420 ;
        RECT 2380.020 -23.430 2383.020 -23.420 ;
        RECT 2560.020 -23.430 2563.020 -23.420 ;
        RECT 2740.020 -23.430 2743.020 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT 130.020 -28.120 133.020 3547.800 ;
        RECT 310.020 -28.120 313.020 3547.800 ;
        RECT 490.020 -28.120 493.020 3547.800 ;
        RECT 670.020 -28.120 673.020 3547.800 ;
        RECT 850.020 -28.120 853.020 3547.800 ;
        RECT 1030.020 -28.120 1033.020 3547.800 ;
        RECT 1210.020 -28.120 1213.020 3547.800 ;
        RECT 1390.020 -28.120 1393.020 3547.800 ;
        RECT 1570.020 -28.120 1573.020 3547.800 ;
        RECT 1750.020 -28.120 1753.020 3547.800 ;
        RECT 1930.020 -28.120 1933.020 3547.800 ;
        RECT 2110.020 -28.120 2113.020 3547.800 ;
        RECT 2290.020 -28.120 2293.020 3547.800 ;
        RECT 2470.020 -28.120 2473.020 3547.800 ;
        RECT 2650.020 -28.120 2653.020 3547.800 ;
        RECT 2830.020 -28.120 2833.020 3547.800 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
      LAYER via4 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT -32.570 3377.090 -31.390 3378.270 ;
        RECT -32.570 3375.490 -31.390 3376.670 ;
        RECT -32.570 3197.090 -31.390 3198.270 ;
        RECT -32.570 3195.490 -31.390 3196.670 ;
        RECT -32.570 3017.090 -31.390 3018.270 ;
        RECT -32.570 3015.490 -31.390 3016.670 ;
        RECT -32.570 2837.090 -31.390 2838.270 ;
        RECT -32.570 2835.490 -31.390 2836.670 ;
        RECT -32.570 2657.090 -31.390 2658.270 ;
        RECT -32.570 2655.490 -31.390 2656.670 ;
        RECT -32.570 2477.090 -31.390 2478.270 ;
        RECT -32.570 2475.490 -31.390 2476.670 ;
        RECT -32.570 2297.090 -31.390 2298.270 ;
        RECT -32.570 2295.490 -31.390 2296.670 ;
        RECT -32.570 2117.090 -31.390 2118.270 ;
        RECT -32.570 2115.490 -31.390 2116.670 ;
        RECT -32.570 1937.090 -31.390 1938.270 ;
        RECT -32.570 1935.490 -31.390 1936.670 ;
        RECT -32.570 1757.090 -31.390 1758.270 ;
        RECT -32.570 1755.490 -31.390 1756.670 ;
        RECT -32.570 1577.090 -31.390 1578.270 ;
        RECT -32.570 1575.490 -31.390 1576.670 ;
        RECT -32.570 1397.090 -31.390 1398.270 ;
        RECT -32.570 1395.490 -31.390 1396.670 ;
        RECT -32.570 1217.090 -31.390 1218.270 ;
        RECT -32.570 1215.490 -31.390 1216.670 ;
        RECT -32.570 1037.090 -31.390 1038.270 ;
        RECT -32.570 1035.490 -31.390 1036.670 ;
        RECT -32.570 857.090 -31.390 858.270 ;
        RECT -32.570 855.490 -31.390 856.670 ;
        RECT -32.570 677.090 -31.390 678.270 ;
        RECT -32.570 675.490 -31.390 676.670 ;
        RECT -32.570 497.090 -31.390 498.270 ;
        RECT -32.570 495.490 -31.390 496.670 ;
        RECT -32.570 317.090 -31.390 318.270 ;
        RECT -32.570 315.490 -31.390 316.670 ;
        RECT -32.570 137.090 -31.390 138.270 ;
        RECT -32.570 135.490 -31.390 136.670 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 130.930 3546.510 132.110 3547.690 ;
        RECT 130.930 3544.910 132.110 3546.090 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -26.410 132.110 -25.230 ;
        RECT 130.930 -28.010 132.110 -26.830 ;
        RECT 310.930 3546.510 312.110 3547.690 ;
        RECT 310.930 3544.910 312.110 3546.090 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 310.930 2657.090 312.110 2658.270 ;
        RECT 310.930 2655.490 312.110 2656.670 ;
        RECT 310.930 2477.090 312.110 2478.270 ;
        RECT 310.930 2475.490 312.110 2476.670 ;
        RECT 310.930 2297.090 312.110 2298.270 ;
        RECT 310.930 2295.490 312.110 2296.670 ;
        RECT 310.930 2117.090 312.110 2118.270 ;
        RECT 310.930 2115.490 312.110 2116.670 ;
        RECT 310.930 1937.090 312.110 1938.270 ;
        RECT 310.930 1935.490 312.110 1936.670 ;
        RECT 310.930 1757.090 312.110 1758.270 ;
        RECT 310.930 1755.490 312.110 1756.670 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -26.410 312.110 -25.230 ;
        RECT 310.930 -28.010 312.110 -26.830 ;
        RECT 490.930 3546.510 492.110 3547.690 ;
        RECT 490.930 3544.910 492.110 3546.090 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 490.930 3197.090 492.110 3198.270 ;
        RECT 490.930 3195.490 492.110 3196.670 ;
        RECT 490.930 3017.090 492.110 3018.270 ;
        RECT 490.930 3015.490 492.110 3016.670 ;
        RECT 490.930 2837.090 492.110 2838.270 ;
        RECT 490.930 2835.490 492.110 2836.670 ;
        RECT 490.930 2657.090 492.110 2658.270 ;
        RECT 490.930 2655.490 492.110 2656.670 ;
        RECT 490.930 2477.090 492.110 2478.270 ;
        RECT 490.930 2475.490 492.110 2476.670 ;
        RECT 490.930 2297.090 492.110 2298.270 ;
        RECT 490.930 2295.490 492.110 2296.670 ;
        RECT 490.930 2117.090 492.110 2118.270 ;
        RECT 490.930 2115.490 492.110 2116.670 ;
        RECT 490.930 1937.090 492.110 1938.270 ;
        RECT 490.930 1935.490 492.110 1936.670 ;
        RECT 490.930 1757.090 492.110 1758.270 ;
        RECT 490.930 1755.490 492.110 1756.670 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -26.410 492.110 -25.230 ;
        RECT 490.930 -28.010 492.110 -26.830 ;
        RECT 670.930 3546.510 672.110 3547.690 ;
        RECT 670.930 3544.910 672.110 3546.090 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 670.930 3197.090 672.110 3198.270 ;
        RECT 670.930 3195.490 672.110 3196.670 ;
        RECT 670.930 3017.090 672.110 3018.270 ;
        RECT 670.930 3015.490 672.110 3016.670 ;
        RECT 670.930 2837.090 672.110 2838.270 ;
        RECT 670.930 2835.490 672.110 2836.670 ;
        RECT 670.930 2657.090 672.110 2658.270 ;
        RECT 670.930 2655.490 672.110 2656.670 ;
        RECT 670.930 2477.090 672.110 2478.270 ;
        RECT 670.930 2475.490 672.110 2476.670 ;
        RECT 670.930 2297.090 672.110 2298.270 ;
        RECT 670.930 2295.490 672.110 2296.670 ;
        RECT 670.930 2117.090 672.110 2118.270 ;
        RECT 670.930 2115.490 672.110 2116.670 ;
        RECT 670.930 1937.090 672.110 1938.270 ;
        RECT 670.930 1935.490 672.110 1936.670 ;
        RECT 670.930 1757.090 672.110 1758.270 ;
        RECT 670.930 1755.490 672.110 1756.670 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 670.930 857.090 672.110 858.270 ;
        RECT 670.930 855.490 672.110 856.670 ;
        RECT 670.930 677.090 672.110 678.270 ;
        RECT 670.930 675.490 672.110 676.670 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -26.410 672.110 -25.230 ;
        RECT 670.930 -28.010 672.110 -26.830 ;
        RECT 850.930 3546.510 852.110 3547.690 ;
        RECT 850.930 3544.910 852.110 3546.090 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 850.930 2657.090 852.110 2658.270 ;
        RECT 850.930 2655.490 852.110 2656.670 ;
        RECT 850.930 2477.090 852.110 2478.270 ;
        RECT 850.930 2475.490 852.110 2476.670 ;
        RECT 850.930 2297.090 852.110 2298.270 ;
        RECT 850.930 2295.490 852.110 2296.670 ;
        RECT 850.930 2117.090 852.110 2118.270 ;
        RECT 850.930 2115.490 852.110 2116.670 ;
        RECT 850.930 1937.090 852.110 1938.270 ;
        RECT 850.930 1935.490 852.110 1936.670 ;
        RECT 850.930 1757.090 852.110 1758.270 ;
        RECT 850.930 1755.490 852.110 1756.670 ;
        RECT 850.930 1577.090 852.110 1578.270 ;
        RECT 850.930 1575.490 852.110 1576.670 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 850.930 857.090 852.110 858.270 ;
        RECT 850.930 855.490 852.110 856.670 ;
        RECT 850.930 677.090 852.110 678.270 ;
        RECT 850.930 675.490 852.110 676.670 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -26.410 852.110 -25.230 ;
        RECT 850.930 -28.010 852.110 -26.830 ;
        RECT 1030.930 3546.510 1032.110 3547.690 ;
        RECT 1030.930 3544.910 1032.110 3546.090 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1030.930 3197.090 1032.110 3198.270 ;
        RECT 1030.930 3195.490 1032.110 3196.670 ;
        RECT 1030.930 3017.090 1032.110 3018.270 ;
        RECT 1030.930 3015.490 1032.110 3016.670 ;
        RECT 1030.930 2837.090 1032.110 2838.270 ;
        RECT 1030.930 2835.490 1032.110 2836.670 ;
        RECT 1030.930 2657.090 1032.110 2658.270 ;
        RECT 1030.930 2655.490 1032.110 2656.670 ;
        RECT 1030.930 2477.090 1032.110 2478.270 ;
        RECT 1030.930 2475.490 1032.110 2476.670 ;
        RECT 1030.930 2297.090 1032.110 2298.270 ;
        RECT 1030.930 2295.490 1032.110 2296.670 ;
        RECT 1030.930 2117.090 1032.110 2118.270 ;
        RECT 1030.930 2115.490 1032.110 2116.670 ;
        RECT 1030.930 1937.090 1032.110 1938.270 ;
        RECT 1030.930 1935.490 1032.110 1936.670 ;
        RECT 1030.930 1757.090 1032.110 1758.270 ;
        RECT 1030.930 1755.490 1032.110 1756.670 ;
        RECT 1030.930 1577.090 1032.110 1578.270 ;
        RECT 1030.930 1575.490 1032.110 1576.670 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1030.930 857.090 1032.110 858.270 ;
        RECT 1030.930 855.490 1032.110 856.670 ;
        RECT 1030.930 677.090 1032.110 678.270 ;
        RECT 1030.930 675.490 1032.110 676.670 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -26.410 1032.110 -25.230 ;
        RECT 1030.930 -28.010 1032.110 -26.830 ;
        RECT 1210.930 3546.510 1212.110 3547.690 ;
        RECT 1210.930 3544.910 1212.110 3546.090 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1210.930 3197.090 1212.110 3198.270 ;
        RECT 1210.930 3195.490 1212.110 3196.670 ;
        RECT 1210.930 3017.090 1212.110 3018.270 ;
        RECT 1210.930 3015.490 1212.110 3016.670 ;
        RECT 1210.930 2837.090 1212.110 2838.270 ;
        RECT 1210.930 2835.490 1212.110 2836.670 ;
        RECT 1210.930 2657.090 1212.110 2658.270 ;
        RECT 1210.930 2655.490 1212.110 2656.670 ;
        RECT 1210.930 2477.090 1212.110 2478.270 ;
        RECT 1210.930 2475.490 1212.110 2476.670 ;
        RECT 1210.930 2297.090 1212.110 2298.270 ;
        RECT 1210.930 2295.490 1212.110 2296.670 ;
        RECT 1210.930 2117.090 1212.110 2118.270 ;
        RECT 1210.930 2115.490 1212.110 2116.670 ;
        RECT 1210.930 1937.090 1212.110 1938.270 ;
        RECT 1210.930 1935.490 1212.110 1936.670 ;
        RECT 1210.930 1757.090 1212.110 1758.270 ;
        RECT 1210.930 1755.490 1212.110 1756.670 ;
        RECT 1210.930 1577.090 1212.110 1578.270 ;
        RECT 1210.930 1575.490 1212.110 1576.670 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1210.930 857.090 1212.110 858.270 ;
        RECT 1210.930 855.490 1212.110 856.670 ;
        RECT 1210.930 677.090 1212.110 678.270 ;
        RECT 1210.930 675.490 1212.110 676.670 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -26.410 1212.110 -25.230 ;
        RECT 1210.930 -28.010 1212.110 -26.830 ;
        RECT 1390.930 3546.510 1392.110 3547.690 ;
        RECT 1390.930 3544.910 1392.110 3546.090 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1390.930 2657.090 1392.110 2658.270 ;
        RECT 1390.930 2655.490 1392.110 2656.670 ;
        RECT 1390.930 2477.090 1392.110 2478.270 ;
        RECT 1390.930 2475.490 1392.110 2476.670 ;
        RECT 1390.930 2297.090 1392.110 2298.270 ;
        RECT 1390.930 2295.490 1392.110 2296.670 ;
        RECT 1390.930 2117.090 1392.110 2118.270 ;
        RECT 1390.930 2115.490 1392.110 2116.670 ;
        RECT 1390.930 1937.090 1392.110 1938.270 ;
        RECT 1390.930 1935.490 1392.110 1936.670 ;
        RECT 1390.930 1757.090 1392.110 1758.270 ;
        RECT 1390.930 1755.490 1392.110 1756.670 ;
        RECT 1390.930 1577.090 1392.110 1578.270 ;
        RECT 1390.930 1575.490 1392.110 1576.670 ;
        RECT 1390.930 1397.090 1392.110 1398.270 ;
        RECT 1390.930 1395.490 1392.110 1396.670 ;
        RECT 1390.930 1217.090 1392.110 1218.270 ;
        RECT 1390.930 1215.490 1392.110 1216.670 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1390.930 857.090 1392.110 858.270 ;
        RECT 1390.930 855.490 1392.110 856.670 ;
        RECT 1390.930 677.090 1392.110 678.270 ;
        RECT 1390.930 675.490 1392.110 676.670 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -26.410 1392.110 -25.230 ;
        RECT 1390.930 -28.010 1392.110 -26.830 ;
        RECT 1570.930 3546.510 1572.110 3547.690 ;
        RECT 1570.930 3544.910 1572.110 3546.090 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1570.930 3017.090 1572.110 3018.270 ;
        RECT 1570.930 3015.490 1572.110 3016.670 ;
        RECT 1570.930 2837.090 1572.110 2838.270 ;
        RECT 1570.930 2835.490 1572.110 2836.670 ;
        RECT 1570.930 2657.090 1572.110 2658.270 ;
        RECT 1570.930 2655.490 1572.110 2656.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1570.930 2297.090 1572.110 2298.270 ;
        RECT 1570.930 2295.490 1572.110 2296.670 ;
        RECT 1570.930 2117.090 1572.110 2118.270 ;
        RECT 1570.930 2115.490 1572.110 2116.670 ;
        RECT 1570.930 1937.090 1572.110 1938.270 ;
        RECT 1570.930 1935.490 1572.110 1936.670 ;
        RECT 1570.930 1757.090 1572.110 1758.270 ;
        RECT 1570.930 1755.490 1572.110 1756.670 ;
        RECT 1570.930 1577.090 1572.110 1578.270 ;
        RECT 1570.930 1575.490 1572.110 1576.670 ;
        RECT 1570.930 1397.090 1572.110 1398.270 ;
        RECT 1570.930 1395.490 1572.110 1396.670 ;
        RECT 1570.930 1217.090 1572.110 1218.270 ;
        RECT 1570.930 1215.490 1572.110 1216.670 ;
        RECT 1570.930 1037.090 1572.110 1038.270 ;
        RECT 1570.930 1035.490 1572.110 1036.670 ;
        RECT 1570.930 857.090 1572.110 858.270 ;
        RECT 1570.930 855.490 1572.110 856.670 ;
        RECT 1570.930 677.090 1572.110 678.270 ;
        RECT 1570.930 675.490 1572.110 676.670 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -26.410 1572.110 -25.230 ;
        RECT 1570.930 -28.010 1572.110 -26.830 ;
        RECT 1750.930 3546.510 1752.110 3547.690 ;
        RECT 1750.930 3544.910 1752.110 3546.090 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1750.930 3017.090 1752.110 3018.270 ;
        RECT 1750.930 3015.490 1752.110 3016.670 ;
        RECT 1750.930 2837.090 1752.110 2838.270 ;
        RECT 1750.930 2835.490 1752.110 2836.670 ;
        RECT 1750.930 2657.090 1752.110 2658.270 ;
        RECT 1750.930 2655.490 1752.110 2656.670 ;
        RECT 1750.930 2477.090 1752.110 2478.270 ;
        RECT 1750.930 2475.490 1752.110 2476.670 ;
        RECT 1750.930 2297.090 1752.110 2298.270 ;
        RECT 1750.930 2295.490 1752.110 2296.670 ;
        RECT 1750.930 2117.090 1752.110 2118.270 ;
        RECT 1750.930 2115.490 1752.110 2116.670 ;
        RECT 1750.930 1937.090 1752.110 1938.270 ;
        RECT 1750.930 1935.490 1752.110 1936.670 ;
        RECT 1750.930 1757.090 1752.110 1758.270 ;
        RECT 1750.930 1755.490 1752.110 1756.670 ;
        RECT 1750.930 1577.090 1752.110 1578.270 ;
        RECT 1750.930 1575.490 1752.110 1576.670 ;
        RECT 1750.930 1397.090 1752.110 1398.270 ;
        RECT 1750.930 1395.490 1752.110 1396.670 ;
        RECT 1750.930 1217.090 1752.110 1218.270 ;
        RECT 1750.930 1215.490 1752.110 1216.670 ;
        RECT 1750.930 1037.090 1752.110 1038.270 ;
        RECT 1750.930 1035.490 1752.110 1036.670 ;
        RECT 1750.930 857.090 1752.110 858.270 ;
        RECT 1750.930 855.490 1752.110 856.670 ;
        RECT 1750.930 677.090 1752.110 678.270 ;
        RECT 1750.930 675.490 1752.110 676.670 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -26.410 1752.110 -25.230 ;
        RECT 1750.930 -28.010 1752.110 -26.830 ;
        RECT 1930.930 3546.510 1932.110 3547.690 ;
        RECT 1930.930 3544.910 1932.110 3546.090 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 1930.930 2837.090 1932.110 2838.270 ;
        RECT 1930.930 2835.490 1932.110 2836.670 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 1930.930 2477.090 1932.110 2478.270 ;
        RECT 1930.930 2475.490 1932.110 2476.670 ;
        RECT 1930.930 2297.090 1932.110 2298.270 ;
        RECT 1930.930 2295.490 1932.110 2296.670 ;
        RECT 1930.930 2117.090 1932.110 2118.270 ;
        RECT 1930.930 2115.490 1932.110 2116.670 ;
        RECT 1930.930 1937.090 1932.110 1938.270 ;
        RECT 1930.930 1935.490 1932.110 1936.670 ;
        RECT 1930.930 1757.090 1932.110 1758.270 ;
        RECT 1930.930 1755.490 1932.110 1756.670 ;
        RECT 1930.930 1577.090 1932.110 1578.270 ;
        RECT 1930.930 1575.490 1932.110 1576.670 ;
        RECT 1930.930 1397.090 1932.110 1398.270 ;
        RECT 1930.930 1395.490 1932.110 1396.670 ;
        RECT 1930.930 1217.090 1932.110 1218.270 ;
        RECT 1930.930 1215.490 1932.110 1216.670 ;
        RECT 1930.930 1037.090 1932.110 1038.270 ;
        RECT 1930.930 1035.490 1932.110 1036.670 ;
        RECT 1930.930 857.090 1932.110 858.270 ;
        RECT 1930.930 855.490 1932.110 856.670 ;
        RECT 1930.930 677.090 1932.110 678.270 ;
        RECT 1930.930 675.490 1932.110 676.670 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -26.410 1932.110 -25.230 ;
        RECT 1930.930 -28.010 1932.110 -26.830 ;
        RECT 2110.930 3546.510 2112.110 3547.690 ;
        RECT 2110.930 3544.910 2112.110 3546.090 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2110.930 2657.090 2112.110 2658.270 ;
        RECT 2110.930 2655.490 2112.110 2656.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2110.930 2297.090 2112.110 2298.270 ;
        RECT 2110.930 2295.490 2112.110 2296.670 ;
        RECT 2110.930 2117.090 2112.110 2118.270 ;
        RECT 2110.930 2115.490 2112.110 2116.670 ;
        RECT 2110.930 1937.090 2112.110 1938.270 ;
        RECT 2110.930 1935.490 2112.110 1936.670 ;
        RECT 2110.930 1757.090 2112.110 1758.270 ;
        RECT 2110.930 1755.490 2112.110 1756.670 ;
        RECT 2110.930 1577.090 2112.110 1578.270 ;
        RECT 2110.930 1575.490 2112.110 1576.670 ;
        RECT 2110.930 1397.090 2112.110 1398.270 ;
        RECT 2110.930 1395.490 2112.110 1396.670 ;
        RECT 2110.930 1217.090 2112.110 1218.270 ;
        RECT 2110.930 1215.490 2112.110 1216.670 ;
        RECT 2110.930 1037.090 2112.110 1038.270 ;
        RECT 2110.930 1035.490 2112.110 1036.670 ;
        RECT 2110.930 857.090 2112.110 858.270 ;
        RECT 2110.930 855.490 2112.110 856.670 ;
        RECT 2110.930 677.090 2112.110 678.270 ;
        RECT 2110.930 675.490 2112.110 676.670 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -26.410 2112.110 -25.230 ;
        RECT 2110.930 -28.010 2112.110 -26.830 ;
        RECT 2290.930 3546.510 2292.110 3547.690 ;
        RECT 2290.930 3544.910 2292.110 3546.090 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2290.930 3017.090 2292.110 3018.270 ;
        RECT 2290.930 3015.490 2292.110 3016.670 ;
        RECT 2290.930 2837.090 2292.110 2838.270 ;
        RECT 2290.930 2835.490 2292.110 2836.670 ;
        RECT 2290.930 2657.090 2292.110 2658.270 ;
        RECT 2290.930 2655.490 2292.110 2656.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2290.930 2297.090 2292.110 2298.270 ;
        RECT 2290.930 2295.490 2292.110 2296.670 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2290.930 1937.090 2292.110 1938.270 ;
        RECT 2290.930 1935.490 2292.110 1936.670 ;
        RECT 2290.930 1757.090 2292.110 1758.270 ;
        RECT 2290.930 1755.490 2292.110 1756.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2290.930 1397.090 2292.110 1398.270 ;
        RECT 2290.930 1395.490 2292.110 1396.670 ;
        RECT 2290.930 1217.090 2292.110 1218.270 ;
        RECT 2290.930 1215.490 2292.110 1216.670 ;
        RECT 2290.930 1037.090 2292.110 1038.270 ;
        RECT 2290.930 1035.490 2292.110 1036.670 ;
        RECT 2290.930 857.090 2292.110 858.270 ;
        RECT 2290.930 855.490 2292.110 856.670 ;
        RECT 2290.930 677.090 2292.110 678.270 ;
        RECT 2290.930 675.490 2292.110 676.670 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -26.410 2292.110 -25.230 ;
        RECT 2290.930 -28.010 2292.110 -26.830 ;
        RECT 2470.930 3546.510 2472.110 3547.690 ;
        RECT 2470.930 3544.910 2472.110 3546.090 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2470.930 3017.090 2472.110 3018.270 ;
        RECT 2470.930 3015.490 2472.110 3016.670 ;
        RECT 2470.930 2837.090 2472.110 2838.270 ;
        RECT 2470.930 2835.490 2472.110 2836.670 ;
        RECT 2470.930 2657.090 2472.110 2658.270 ;
        RECT 2470.930 2655.490 2472.110 2656.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2470.930 2297.090 2472.110 2298.270 ;
        RECT 2470.930 2295.490 2472.110 2296.670 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2470.930 1937.090 2472.110 1938.270 ;
        RECT 2470.930 1935.490 2472.110 1936.670 ;
        RECT 2470.930 1757.090 2472.110 1758.270 ;
        RECT 2470.930 1755.490 2472.110 1756.670 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2470.930 1397.090 2472.110 1398.270 ;
        RECT 2470.930 1395.490 2472.110 1396.670 ;
        RECT 2470.930 1217.090 2472.110 1218.270 ;
        RECT 2470.930 1215.490 2472.110 1216.670 ;
        RECT 2470.930 1037.090 2472.110 1038.270 ;
        RECT 2470.930 1035.490 2472.110 1036.670 ;
        RECT 2470.930 857.090 2472.110 858.270 ;
        RECT 2470.930 855.490 2472.110 856.670 ;
        RECT 2470.930 677.090 2472.110 678.270 ;
        RECT 2470.930 675.490 2472.110 676.670 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -26.410 2472.110 -25.230 ;
        RECT 2470.930 -28.010 2472.110 -26.830 ;
        RECT 2650.930 3546.510 2652.110 3547.690 ;
        RECT 2650.930 3544.910 2652.110 3546.090 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -26.410 2652.110 -25.230 ;
        RECT 2650.930 -28.010 2652.110 -26.830 ;
        RECT 2830.930 3546.510 2832.110 3547.690 ;
        RECT 2830.930 3544.910 2832.110 3546.090 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -26.410 2832.110 -25.230 ;
        RECT 2830.930 -28.010 2832.110 -26.830 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT 2951.010 3377.090 2952.190 3378.270 ;
        RECT 2951.010 3375.490 2952.190 3376.670 ;
        RECT 2951.010 3197.090 2952.190 3198.270 ;
        RECT 2951.010 3195.490 2952.190 3196.670 ;
        RECT 2951.010 3017.090 2952.190 3018.270 ;
        RECT 2951.010 3015.490 2952.190 3016.670 ;
        RECT 2951.010 2837.090 2952.190 2838.270 ;
        RECT 2951.010 2835.490 2952.190 2836.670 ;
        RECT 2951.010 2657.090 2952.190 2658.270 ;
        RECT 2951.010 2655.490 2952.190 2656.670 ;
        RECT 2951.010 2477.090 2952.190 2478.270 ;
        RECT 2951.010 2475.490 2952.190 2476.670 ;
        RECT 2951.010 2297.090 2952.190 2298.270 ;
        RECT 2951.010 2295.490 2952.190 2296.670 ;
        RECT 2951.010 2117.090 2952.190 2118.270 ;
        RECT 2951.010 2115.490 2952.190 2116.670 ;
        RECT 2951.010 1937.090 2952.190 1938.270 ;
        RECT 2951.010 1935.490 2952.190 1936.670 ;
        RECT 2951.010 1757.090 2952.190 1758.270 ;
        RECT 2951.010 1755.490 2952.190 1756.670 ;
        RECT 2951.010 1577.090 2952.190 1578.270 ;
        RECT 2951.010 1575.490 2952.190 1576.670 ;
        RECT 2951.010 1397.090 2952.190 1398.270 ;
        RECT 2951.010 1395.490 2952.190 1396.670 ;
        RECT 2951.010 1217.090 2952.190 1218.270 ;
        RECT 2951.010 1215.490 2952.190 1216.670 ;
        RECT 2951.010 1037.090 2952.190 1038.270 ;
        RECT 2951.010 1035.490 2952.190 1036.670 ;
        RECT 2951.010 857.090 2952.190 858.270 ;
        RECT 2951.010 855.490 2952.190 856.670 ;
        RECT 2951.010 677.090 2952.190 678.270 ;
        RECT 2951.010 675.490 2952.190 676.670 ;
        RECT 2951.010 497.090 2952.190 498.270 ;
        RECT 2951.010 495.490 2952.190 496.670 ;
        RECT 2951.010 317.090 2952.190 318.270 ;
        RECT 2951.010 315.490 2952.190 316.670 ;
        RECT 2951.010 137.090 2952.190 138.270 ;
        RECT 2951.010 135.490 2952.190 136.670 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
      LAYER met5 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 130.020 3547.800 133.020 3547.810 ;
        RECT 310.020 3547.800 313.020 3547.810 ;
        RECT 490.020 3547.800 493.020 3547.810 ;
        RECT 670.020 3547.800 673.020 3547.810 ;
        RECT 850.020 3547.800 853.020 3547.810 ;
        RECT 1030.020 3547.800 1033.020 3547.810 ;
        RECT 1210.020 3547.800 1213.020 3547.810 ;
        RECT 1390.020 3547.800 1393.020 3547.810 ;
        RECT 1570.020 3547.800 1573.020 3547.810 ;
        RECT 1750.020 3547.800 1753.020 3547.810 ;
        RECT 1930.020 3547.800 1933.020 3547.810 ;
        RECT 2110.020 3547.800 2113.020 3547.810 ;
        RECT 2290.020 3547.800 2293.020 3547.810 ;
        RECT 2470.020 3547.800 2473.020 3547.810 ;
        RECT 2650.020 3547.800 2653.020 3547.810 ;
        RECT 2830.020 3547.800 2833.020 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 130.020 3544.790 133.020 3544.800 ;
        RECT 310.020 3544.790 313.020 3544.800 ;
        RECT 490.020 3544.790 493.020 3544.800 ;
        RECT 670.020 3544.790 673.020 3544.800 ;
        RECT 850.020 3544.790 853.020 3544.800 ;
        RECT 1030.020 3544.790 1033.020 3544.800 ;
        RECT 1210.020 3544.790 1213.020 3544.800 ;
        RECT 1390.020 3544.790 1393.020 3544.800 ;
        RECT 1570.020 3544.790 1573.020 3544.800 ;
        RECT 1750.020 3544.790 1753.020 3544.800 ;
        RECT 1930.020 3544.790 1933.020 3544.800 ;
        RECT 2110.020 3544.790 2113.020 3544.800 ;
        RECT 2290.020 3544.790 2293.020 3544.800 ;
        RECT 2470.020 3544.790 2473.020 3544.800 ;
        RECT 2650.020 3544.790 2653.020 3544.800 ;
        RECT 2830.020 3544.790 2833.020 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -33.480 3378.380 -30.480 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2950.100 3378.380 2953.100 3378.390 ;
        RECT -33.480 3375.380 2953.100 3378.380 ;
        RECT -33.480 3375.370 -30.480 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2950.100 3375.370 2953.100 3375.380 ;
        RECT -33.480 3198.380 -30.480 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 490.020 3198.380 493.020 3198.390 ;
        RECT 670.020 3198.380 673.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1030.020 3198.380 1033.020 3198.390 ;
        RECT 1210.020 3198.380 1213.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2950.100 3198.380 2953.100 3198.390 ;
        RECT -33.480 3195.380 2953.100 3198.380 ;
        RECT -33.480 3195.370 -30.480 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 490.020 3195.370 493.020 3195.380 ;
        RECT 670.020 3195.370 673.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1030.020 3195.370 1033.020 3195.380 ;
        RECT 1210.020 3195.370 1213.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2950.100 3195.370 2953.100 3195.380 ;
        RECT -33.480 3018.380 -30.480 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 490.020 3018.380 493.020 3018.390 ;
        RECT 670.020 3018.380 673.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1030.020 3018.380 1033.020 3018.390 ;
        RECT 1210.020 3018.380 1213.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1570.020 3018.380 1573.020 3018.390 ;
        RECT 1750.020 3018.380 1753.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2290.020 3018.380 2293.020 3018.390 ;
        RECT 2470.020 3018.380 2473.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2950.100 3018.380 2953.100 3018.390 ;
        RECT -33.480 3015.380 2953.100 3018.380 ;
        RECT -33.480 3015.370 -30.480 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 490.020 3015.370 493.020 3015.380 ;
        RECT 670.020 3015.370 673.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1030.020 3015.370 1033.020 3015.380 ;
        RECT 1210.020 3015.370 1213.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1570.020 3015.370 1573.020 3015.380 ;
        RECT 1750.020 3015.370 1753.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2290.020 3015.370 2293.020 3015.380 ;
        RECT 2470.020 3015.370 2473.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2950.100 3015.370 2953.100 3015.380 ;
        RECT -33.480 2838.380 -30.480 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 490.020 2838.380 493.020 2838.390 ;
        RECT 670.020 2838.380 673.020 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1030.020 2838.380 1033.020 2838.390 ;
        RECT 1210.020 2838.380 1213.020 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1570.020 2838.380 1573.020 2838.390 ;
        RECT 1750.020 2838.380 1753.020 2838.390 ;
        RECT 1930.020 2838.380 1933.020 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2290.020 2838.380 2293.020 2838.390 ;
        RECT 2470.020 2838.380 2473.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2950.100 2838.380 2953.100 2838.390 ;
        RECT -33.480 2835.380 2953.100 2838.380 ;
        RECT -33.480 2835.370 -30.480 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 490.020 2835.370 493.020 2835.380 ;
        RECT 670.020 2835.370 673.020 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1030.020 2835.370 1033.020 2835.380 ;
        RECT 1210.020 2835.370 1213.020 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1570.020 2835.370 1573.020 2835.380 ;
        RECT 1750.020 2835.370 1753.020 2835.380 ;
        RECT 1930.020 2835.370 1933.020 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2290.020 2835.370 2293.020 2835.380 ;
        RECT 2470.020 2835.370 2473.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2950.100 2835.370 2953.100 2835.380 ;
        RECT -33.480 2658.380 -30.480 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 310.020 2658.380 313.020 2658.390 ;
        RECT 490.020 2658.380 493.020 2658.390 ;
        RECT 670.020 2658.380 673.020 2658.390 ;
        RECT 850.020 2658.380 853.020 2658.390 ;
        RECT 1030.020 2658.380 1033.020 2658.390 ;
        RECT 1210.020 2658.380 1213.020 2658.390 ;
        RECT 1390.020 2658.380 1393.020 2658.390 ;
        RECT 1570.020 2658.380 1573.020 2658.390 ;
        RECT 1750.020 2658.380 1753.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2110.020 2658.380 2113.020 2658.390 ;
        RECT 2290.020 2658.380 2293.020 2658.390 ;
        RECT 2470.020 2658.380 2473.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2950.100 2658.380 2953.100 2658.390 ;
        RECT -33.480 2655.380 2953.100 2658.380 ;
        RECT -33.480 2655.370 -30.480 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 310.020 2655.370 313.020 2655.380 ;
        RECT 490.020 2655.370 493.020 2655.380 ;
        RECT 670.020 2655.370 673.020 2655.380 ;
        RECT 850.020 2655.370 853.020 2655.380 ;
        RECT 1030.020 2655.370 1033.020 2655.380 ;
        RECT 1210.020 2655.370 1213.020 2655.380 ;
        RECT 1390.020 2655.370 1393.020 2655.380 ;
        RECT 1570.020 2655.370 1573.020 2655.380 ;
        RECT 1750.020 2655.370 1753.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2110.020 2655.370 2113.020 2655.380 ;
        RECT 2290.020 2655.370 2293.020 2655.380 ;
        RECT 2470.020 2655.370 2473.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2950.100 2655.370 2953.100 2655.380 ;
        RECT -33.480 2478.380 -30.480 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 310.020 2478.380 313.020 2478.390 ;
        RECT 490.020 2478.380 493.020 2478.390 ;
        RECT 670.020 2478.380 673.020 2478.390 ;
        RECT 850.020 2478.380 853.020 2478.390 ;
        RECT 1030.020 2478.380 1033.020 2478.390 ;
        RECT 1210.020 2478.380 1213.020 2478.390 ;
        RECT 1390.020 2478.380 1393.020 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 1750.020 2478.380 1753.020 2478.390 ;
        RECT 1930.020 2478.380 1933.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2950.100 2478.380 2953.100 2478.390 ;
        RECT -33.480 2475.380 2953.100 2478.380 ;
        RECT -33.480 2475.370 -30.480 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 310.020 2475.370 313.020 2475.380 ;
        RECT 490.020 2475.370 493.020 2475.380 ;
        RECT 670.020 2475.370 673.020 2475.380 ;
        RECT 850.020 2475.370 853.020 2475.380 ;
        RECT 1030.020 2475.370 1033.020 2475.380 ;
        RECT 1210.020 2475.370 1213.020 2475.380 ;
        RECT 1390.020 2475.370 1393.020 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 1750.020 2475.370 1753.020 2475.380 ;
        RECT 1930.020 2475.370 1933.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2950.100 2475.370 2953.100 2475.380 ;
        RECT -33.480 2298.380 -30.480 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 310.020 2298.380 313.020 2298.390 ;
        RECT 490.020 2298.380 493.020 2298.390 ;
        RECT 670.020 2298.380 673.020 2298.390 ;
        RECT 850.020 2298.380 853.020 2298.390 ;
        RECT 1030.020 2298.380 1033.020 2298.390 ;
        RECT 1210.020 2298.380 1213.020 2298.390 ;
        RECT 1390.020 2298.380 1393.020 2298.390 ;
        RECT 1570.020 2298.380 1573.020 2298.390 ;
        RECT 1750.020 2298.380 1753.020 2298.390 ;
        RECT 1930.020 2298.380 1933.020 2298.390 ;
        RECT 2110.020 2298.380 2113.020 2298.390 ;
        RECT 2290.020 2298.380 2293.020 2298.390 ;
        RECT 2470.020 2298.380 2473.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2950.100 2298.380 2953.100 2298.390 ;
        RECT -33.480 2295.380 2953.100 2298.380 ;
        RECT -33.480 2295.370 -30.480 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 310.020 2295.370 313.020 2295.380 ;
        RECT 490.020 2295.370 493.020 2295.380 ;
        RECT 670.020 2295.370 673.020 2295.380 ;
        RECT 850.020 2295.370 853.020 2295.380 ;
        RECT 1030.020 2295.370 1033.020 2295.380 ;
        RECT 1210.020 2295.370 1213.020 2295.380 ;
        RECT 1390.020 2295.370 1393.020 2295.380 ;
        RECT 1570.020 2295.370 1573.020 2295.380 ;
        RECT 1750.020 2295.370 1753.020 2295.380 ;
        RECT 1930.020 2295.370 1933.020 2295.380 ;
        RECT 2110.020 2295.370 2113.020 2295.380 ;
        RECT 2290.020 2295.370 2293.020 2295.380 ;
        RECT 2470.020 2295.370 2473.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2950.100 2295.370 2953.100 2295.380 ;
        RECT -33.480 2118.380 -30.480 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 310.020 2118.380 313.020 2118.390 ;
        RECT 490.020 2118.380 493.020 2118.390 ;
        RECT 670.020 2118.380 673.020 2118.390 ;
        RECT 850.020 2118.380 853.020 2118.390 ;
        RECT 1030.020 2118.380 1033.020 2118.390 ;
        RECT 1210.020 2118.380 1213.020 2118.390 ;
        RECT 1390.020 2118.380 1393.020 2118.390 ;
        RECT 1570.020 2118.380 1573.020 2118.390 ;
        RECT 1750.020 2118.380 1753.020 2118.390 ;
        RECT 1930.020 2118.380 1933.020 2118.390 ;
        RECT 2110.020 2118.380 2113.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2950.100 2118.380 2953.100 2118.390 ;
        RECT -33.480 2115.380 2953.100 2118.380 ;
        RECT -33.480 2115.370 -30.480 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 310.020 2115.370 313.020 2115.380 ;
        RECT 490.020 2115.370 493.020 2115.380 ;
        RECT 670.020 2115.370 673.020 2115.380 ;
        RECT 850.020 2115.370 853.020 2115.380 ;
        RECT 1030.020 2115.370 1033.020 2115.380 ;
        RECT 1210.020 2115.370 1213.020 2115.380 ;
        RECT 1390.020 2115.370 1393.020 2115.380 ;
        RECT 1570.020 2115.370 1573.020 2115.380 ;
        RECT 1750.020 2115.370 1753.020 2115.380 ;
        RECT 1930.020 2115.370 1933.020 2115.380 ;
        RECT 2110.020 2115.370 2113.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2950.100 2115.370 2953.100 2115.380 ;
        RECT -33.480 1938.380 -30.480 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 310.020 1938.380 313.020 1938.390 ;
        RECT 490.020 1938.380 493.020 1938.390 ;
        RECT 670.020 1938.380 673.020 1938.390 ;
        RECT 850.020 1938.380 853.020 1938.390 ;
        RECT 1030.020 1938.380 1033.020 1938.390 ;
        RECT 1210.020 1938.380 1213.020 1938.390 ;
        RECT 1390.020 1938.380 1393.020 1938.390 ;
        RECT 1570.020 1938.380 1573.020 1938.390 ;
        RECT 1750.020 1938.380 1753.020 1938.390 ;
        RECT 1930.020 1938.380 1933.020 1938.390 ;
        RECT 2110.020 1938.380 2113.020 1938.390 ;
        RECT 2290.020 1938.380 2293.020 1938.390 ;
        RECT 2470.020 1938.380 2473.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2950.100 1938.380 2953.100 1938.390 ;
        RECT -33.480 1935.380 2953.100 1938.380 ;
        RECT -33.480 1935.370 -30.480 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 310.020 1935.370 313.020 1935.380 ;
        RECT 490.020 1935.370 493.020 1935.380 ;
        RECT 670.020 1935.370 673.020 1935.380 ;
        RECT 850.020 1935.370 853.020 1935.380 ;
        RECT 1030.020 1935.370 1033.020 1935.380 ;
        RECT 1210.020 1935.370 1213.020 1935.380 ;
        RECT 1390.020 1935.370 1393.020 1935.380 ;
        RECT 1570.020 1935.370 1573.020 1935.380 ;
        RECT 1750.020 1935.370 1753.020 1935.380 ;
        RECT 1930.020 1935.370 1933.020 1935.380 ;
        RECT 2110.020 1935.370 2113.020 1935.380 ;
        RECT 2290.020 1935.370 2293.020 1935.380 ;
        RECT 2470.020 1935.370 2473.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2950.100 1935.370 2953.100 1935.380 ;
        RECT -33.480 1758.380 -30.480 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 310.020 1758.380 313.020 1758.390 ;
        RECT 490.020 1758.380 493.020 1758.390 ;
        RECT 670.020 1758.380 673.020 1758.390 ;
        RECT 850.020 1758.380 853.020 1758.390 ;
        RECT 1030.020 1758.380 1033.020 1758.390 ;
        RECT 1210.020 1758.380 1213.020 1758.390 ;
        RECT 1390.020 1758.380 1393.020 1758.390 ;
        RECT 1570.020 1758.380 1573.020 1758.390 ;
        RECT 1750.020 1758.380 1753.020 1758.390 ;
        RECT 1930.020 1758.380 1933.020 1758.390 ;
        RECT 2110.020 1758.380 2113.020 1758.390 ;
        RECT 2290.020 1758.380 2293.020 1758.390 ;
        RECT 2470.020 1758.380 2473.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2950.100 1758.380 2953.100 1758.390 ;
        RECT -33.480 1755.380 2953.100 1758.380 ;
        RECT -33.480 1755.370 -30.480 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 310.020 1755.370 313.020 1755.380 ;
        RECT 490.020 1755.370 493.020 1755.380 ;
        RECT 670.020 1755.370 673.020 1755.380 ;
        RECT 850.020 1755.370 853.020 1755.380 ;
        RECT 1030.020 1755.370 1033.020 1755.380 ;
        RECT 1210.020 1755.370 1213.020 1755.380 ;
        RECT 1390.020 1755.370 1393.020 1755.380 ;
        RECT 1570.020 1755.370 1573.020 1755.380 ;
        RECT 1750.020 1755.370 1753.020 1755.380 ;
        RECT 1930.020 1755.370 1933.020 1755.380 ;
        RECT 2110.020 1755.370 2113.020 1755.380 ;
        RECT 2290.020 1755.370 2293.020 1755.380 ;
        RECT 2470.020 1755.370 2473.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2950.100 1755.370 2953.100 1755.380 ;
        RECT -33.480 1578.380 -30.480 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 850.020 1578.380 853.020 1578.390 ;
        RECT 1030.020 1578.380 1033.020 1578.390 ;
        RECT 1210.020 1578.380 1213.020 1578.390 ;
        RECT 1390.020 1578.380 1393.020 1578.390 ;
        RECT 1570.020 1578.380 1573.020 1578.390 ;
        RECT 1750.020 1578.380 1753.020 1578.390 ;
        RECT 1930.020 1578.380 1933.020 1578.390 ;
        RECT 2110.020 1578.380 2113.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2950.100 1578.380 2953.100 1578.390 ;
        RECT -33.480 1575.380 2953.100 1578.380 ;
        RECT -33.480 1575.370 -30.480 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 850.020 1575.370 853.020 1575.380 ;
        RECT 1030.020 1575.370 1033.020 1575.380 ;
        RECT 1210.020 1575.370 1213.020 1575.380 ;
        RECT 1390.020 1575.370 1393.020 1575.380 ;
        RECT 1570.020 1575.370 1573.020 1575.380 ;
        RECT 1750.020 1575.370 1753.020 1575.380 ;
        RECT 1930.020 1575.370 1933.020 1575.380 ;
        RECT 2110.020 1575.370 2113.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2950.100 1575.370 2953.100 1575.380 ;
        RECT -33.480 1398.380 -30.480 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 1390.020 1398.380 1393.020 1398.390 ;
        RECT 1570.020 1398.380 1573.020 1398.390 ;
        RECT 1750.020 1398.380 1753.020 1398.390 ;
        RECT 1930.020 1398.380 1933.020 1398.390 ;
        RECT 2110.020 1398.380 2113.020 1398.390 ;
        RECT 2290.020 1398.380 2293.020 1398.390 ;
        RECT 2470.020 1398.380 2473.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2950.100 1398.380 2953.100 1398.390 ;
        RECT -33.480 1395.380 2953.100 1398.380 ;
        RECT -33.480 1395.370 -30.480 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 1390.020 1395.370 1393.020 1395.380 ;
        RECT 1570.020 1395.370 1573.020 1395.380 ;
        RECT 1750.020 1395.370 1753.020 1395.380 ;
        RECT 1930.020 1395.370 1933.020 1395.380 ;
        RECT 2110.020 1395.370 2113.020 1395.380 ;
        RECT 2290.020 1395.370 2293.020 1395.380 ;
        RECT 2470.020 1395.370 2473.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2950.100 1395.370 2953.100 1395.380 ;
        RECT -33.480 1218.380 -30.480 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 1390.020 1218.380 1393.020 1218.390 ;
        RECT 1570.020 1218.380 1573.020 1218.390 ;
        RECT 1750.020 1218.380 1753.020 1218.390 ;
        RECT 1930.020 1218.380 1933.020 1218.390 ;
        RECT 2110.020 1218.380 2113.020 1218.390 ;
        RECT 2290.020 1218.380 2293.020 1218.390 ;
        RECT 2470.020 1218.380 2473.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2950.100 1218.380 2953.100 1218.390 ;
        RECT -33.480 1215.380 2953.100 1218.380 ;
        RECT -33.480 1215.370 -30.480 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 1390.020 1215.370 1393.020 1215.380 ;
        RECT 1570.020 1215.370 1573.020 1215.380 ;
        RECT 1750.020 1215.370 1753.020 1215.380 ;
        RECT 1930.020 1215.370 1933.020 1215.380 ;
        RECT 2110.020 1215.370 2113.020 1215.380 ;
        RECT 2290.020 1215.370 2293.020 1215.380 ;
        RECT 2470.020 1215.370 2473.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2950.100 1215.370 2953.100 1215.380 ;
        RECT -33.480 1038.380 -30.480 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1570.020 1038.380 1573.020 1038.390 ;
        RECT 1750.020 1038.380 1753.020 1038.390 ;
        RECT 1930.020 1038.380 1933.020 1038.390 ;
        RECT 2110.020 1038.380 2113.020 1038.390 ;
        RECT 2290.020 1038.380 2293.020 1038.390 ;
        RECT 2470.020 1038.380 2473.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2950.100 1038.380 2953.100 1038.390 ;
        RECT -33.480 1035.380 2953.100 1038.380 ;
        RECT -33.480 1035.370 -30.480 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1570.020 1035.370 1573.020 1035.380 ;
        RECT 1750.020 1035.370 1753.020 1035.380 ;
        RECT 1930.020 1035.370 1933.020 1035.380 ;
        RECT 2110.020 1035.370 2113.020 1035.380 ;
        RECT 2290.020 1035.370 2293.020 1035.380 ;
        RECT 2470.020 1035.370 2473.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2950.100 1035.370 2953.100 1035.380 ;
        RECT -33.480 858.380 -30.480 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 670.020 858.380 673.020 858.390 ;
        RECT 850.020 858.380 853.020 858.390 ;
        RECT 1030.020 858.380 1033.020 858.390 ;
        RECT 1210.020 858.380 1213.020 858.390 ;
        RECT 1390.020 858.380 1393.020 858.390 ;
        RECT 1570.020 858.380 1573.020 858.390 ;
        RECT 1750.020 858.380 1753.020 858.390 ;
        RECT 1930.020 858.380 1933.020 858.390 ;
        RECT 2110.020 858.380 2113.020 858.390 ;
        RECT 2290.020 858.380 2293.020 858.390 ;
        RECT 2470.020 858.380 2473.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2950.100 858.380 2953.100 858.390 ;
        RECT -33.480 855.380 2953.100 858.380 ;
        RECT -33.480 855.370 -30.480 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 670.020 855.370 673.020 855.380 ;
        RECT 850.020 855.370 853.020 855.380 ;
        RECT 1030.020 855.370 1033.020 855.380 ;
        RECT 1210.020 855.370 1213.020 855.380 ;
        RECT 1390.020 855.370 1393.020 855.380 ;
        RECT 1570.020 855.370 1573.020 855.380 ;
        RECT 1750.020 855.370 1753.020 855.380 ;
        RECT 1930.020 855.370 1933.020 855.380 ;
        RECT 2110.020 855.370 2113.020 855.380 ;
        RECT 2290.020 855.370 2293.020 855.380 ;
        RECT 2470.020 855.370 2473.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2950.100 855.370 2953.100 855.380 ;
        RECT -33.480 678.380 -30.480 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 670.020 678.380 673.020 678.390 ;
        RECT 850.020 678.380 853.020 678.390 ;
        RECT 1030.020 678.380 1033.020 678.390 ;
        RECT 1210.020 678.380 1213.020 678.390 ;
        RECT 1390.020 678.380 1393.020 678.390 ;
        RECT 1570.020 678.380 1573.020 678.390 ;
        RECT 1750.020 678.380 1753.020 678.390 ;
        RECT 1930.020 678.380 1933.020 678.390 ;
        RECT 2110.020 678.380 2113.020 678.390 ;
        RECT 2290.020 678.380 2293.020 678.390 ;
        RECT 2470.020 678.380 2473.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2950.100 678.380 2953.100 678.390 ;
        RECT -33.480 675.380 2953.100 678.380 ;
        RECT -33.480 675.370 -30.480 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 670.020 675.370 673.020 675.380 ;
        RECT 850.020 675.370 853.020 675.380 ;
        RECT 1030.020 675.370 1033.020 675.380 ;
        RECT 1210.020 675.370 1213.020 675.380 ;
        RECT 1390.020 675.370 1393.020 675.380 ;
        RECT 1570.020 675.370 1573.020 675.380 ;
        RECT 1750.020 675.370 1753.020 675.380 ;
        RECT 1930.020 675.370 1933.020 675.380 ;
        RECT 2110.020 675.370 2113.020 675.380 ;
        RECT 2290.020 675.370 2293.020 675.380 ;
        RECT 2470.020 675.370 2473.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2950.100 675.370 2953.100 675.380 ;
        RECT -33.480 498.380 -30.480 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2950.100 498.380 2953.100 498.390 ;
        RECT -33.480 495.380 2953.100 498.380 ;
        RECT -33.480 495.370 -30.480 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2950.100 495.370 2953.100 495.380 ;
        RECT -33.480 318.380 -30.480 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2950.100 318.380 2953.100 318.390 ;
        RECT -33.480 315.380 2953.100 318.380 ;
        RECT -33.480 315.370 -30.480 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2950.100 315.370 2953.100 315.380 ;
        RECT -33.480 138.380 -30.480 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2950.100 138.380 2953.100 138.390 ;
        RECT -33.480 135.380 2953.100 138.380 ;
        RECT -33.480 135.370 -30.480 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2950.100 135.370 2953.100 135.380 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 130.020 -25.120 133.020 -25.110 ;
        RECT 310.020 -25.120 313.020 -25.110 ;
        RECT 490.020 -25.120 493.020 -25.110 ;
        RECT 670.020 -25.120 673.020 -25.110 ;
        RECT 850.020 -25.120 853.020 -25.110 ;
        RECT 1030.020 -25.120 1033.020 -25.110 ;
        RECT 1210.020 -25.120 1213.020 -25.110 ;
        RECT 1390.020 -25.120 1393.020 -25.110 ;
        RECT 1570.020 -25.120 1573.020 -25.110 ;
        RECT 1750.020 -25.120 1753.020 -25.110 ;
        RECT 1930.020 -25.120 1933.020 -25.110 ;
        RECT 2110.020 -25.120 2113.020 -25.110 ;
        RECT 2290.020 -25.120 2293.020 -25.110 ;
        RECT 2470.020 -25.120 2473.020 -25.110 ;
        RECT 2650.020 -25.120 2653.020 -25.110 ;
        RECT 2830.020 -25.120 2833.020 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 130.020 -28.130 133.020 -28.120 ;
        RECT 310.020 -28.130 313.020 -28.120 ;
        RECT 490.020 -28.130 493.020 -28.120 ;
        RECT 670.020 -28.130 673.020 -28.120 ;
        RECT 850.020 -28.130 853.020 -28.120 ;
        RECT 1030.020 -28.130 1033.020 -28.120 ;
        RECT 1210.020 -28.130 1213.020 -28.120 ;
        RECT 1390.020 -28.130 1393.020 -28.120 ;
        RECT 1570.020 -28.130 1573.020 -28.120 ;
        RECT 1750.020 -28.130 1753.020 -28.120 ;
        RECT 1930.020 -28.130 1933.020 -28.120 ;
        RECT 2110.020 -28.130 2113.020 -28.120 ;
        RECT 2290.020 -28.130 2293.020 -28.120 ;
        RECT 2470.020 -28.130 2473.020 -28.120 ;
        RECT 2650.020 -28.130 2653.020 -28.120 ;
        RECT 2830.020 -28.130 2833.020 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT 58.020 -37.520 61.020 3557.200 ;
        RECT 238.020 -37.520 241.020 3557.200 ;
        RECT 418.020 -37.520 421.020 3557.200 ;
        RECT 598.020 -37.520 601.020 3557.200 ;
        RECT 778.020 -37.520 781.020 3557.200 ;
        RECT 958.020 -37.520 961.020 3557.200 ;
        RECT 1138.020 -37.520 1141.020 3557.200 ;
        RECT 1318.020 -37.520 1321.020 3557.200 ;
        RECT 1498.020 -37.520 1501.020 3557.200 ;
        RECT 1678.020 -37.520 1681.020 3557.200 ;
        RECT 1858.020 -37.520 1861.020 3557.200 ;
        RECT 2038.020 -37.520 2041.020 3557.200 ;
        RECT 2218.020 -37.520 2221.020 3557.200 ;
        RECT 2398.020 -37.520 2401.020 3557.200 ;
        RECT 2578.020 -37.520 2581.020 3557.200 ;
        RECT 2758.020 -37.520 2761.020 3557.200 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT -37.270 3485.090 -36.090 3486.270 ;
        RECT -37.270 3483.490 -36.090 3484.670 ;
        RECT -37.270 3305.090 -36.090 3306.270 ;
        RECT -37.270 3303.490 -36.090 3304.670 ;
        RECT -37.270 3125.090 -36.090 3126.270 ;
        RECT -37.270 3123.490 -36.090 3124.670 ;
        RECT -37.270 2945.090 -36.090 2946.270 ;
        RECT -37.270 2943.490 -36.090 2944.670 ;
        RECT -37.270 2765.090 -36.090 2766.270 ;
        RECT -37.270 2763.490 -36.090 2764.670 ;
        RECT -37.270 2585.090 -36.090 2586.270 ;
        RECT -37.270 2583.490 -36.090 2584.670 ;
        RECT -37.270 2405.090 -36.090 2406.270 ;
        RECT -37.270 2403.490 -36.090 2404.670 ;
        RECT -37.270 2225.090 -36.090 2226.270 ;
        RECT -37.270 2223.490 -36.090 2224.670 ;
        RECT -37.270 2045.090 -36.090 2046.270 ;
        RECT -37.270 2043.490 -36.090 2044.670 ;
        RECT -37.270 1865.090 -36.090 1866.270 ;
        RECT -37.270 1863.490 -36.090 1864.670 ;
        RECT -37.270 1685.090 -36.090 1686.270 ;
        RECT -37.270 1683.490 -36.090 1684.670 ;
        RECT -37.270 1505.090 -36.090 1506.270 ;
        RECT -37.270 1503.490 -36.090 1504.670 ;
        RECT -37.270 1325.090 -36.090 1326.270 ;
        RECT -37.270 1323.490 -36.090 1324.670 ;
        RECT -37.270 1145.090 -36.090 1146.270 ;
        RECT -37.270 1143.490 -36.090 1144.670 ;
        RECT -37.270 965.090 -36.090 966.270 ;
        RECT -37.270 963.490 -36.090 964.670 ;
        RECT -37.270 785.090 -36.090 786.270 ;
        RECT -37.270 783.490 -36.090 784.670 ;
        RECT -37.270 605.090 -36.090 606.270 ;
        RECT -37.270 603.490 -36.090 604.670 ;
        RECT -37.270 425.090 -36.090 426.270 ;
        RECT -37.270 423.490 -36.090 424.670 ;
        RECT -37.270 245.090 -36.090 246.270 ;
        RECT -37.270 243.490 -36.090 244.670 ;
        RECT -37.270 65.090 -36.090 66.270 ;
        RECT -37.270 63.490 -36.090 64.670 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 58.930 3551.210 60.110 3552.390 ;
        RECT 58.930 3549.610 60.110 3550.790 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -31.110 60.110 -29.930 ;
        RECT 58.930 -32.710 60.110 -31.530 ;
        RECT 238.930 3551.210 240.110 3552.390 ;
        RECT 238.930 3549.610 240.110 3550.790 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -31.110 240.110 -29.930 ;
        RECT 238.930 -32.710 240.110 -31.530 ;
        RECT 418.930 3551.210 420.110 3552.390 ;
        RECT 418.930 3549.610 420.110 3550.790 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 418.930 3125.090 420.110 3126.270 ;
        RECT 418.930 3123.490 420.110 3124.670 ;
        RECT 418.930 2945.090 420.110 2946.270 ;
        RECT 418.930 2943.490 420.110 2944.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 418.930 2585.090 420.110 2586.270 ;
        RECT 418.930 2583.490 420.110 2584.670 ;
        RECT 418.930 2405.090 420.110 2406.270 ;
        RECT 418.930 2403.490 420.110 2404.670 ;
        RECT 418.930 2225.090 420.110 2226.270 ;
        RECT 418.930 2223.490 420.110 2224.670 ;
        RECT 418.930 2045.090 420.110 2046.270 ;
        RECT 418.930 2043.490 420.110 2044.670 ;
        RECT 418.930 1865.090 420.110 1866.270 ;
        RECT 418.930 1863.490 420.110 1864.670 ;
        RECT 418.930 1685.090 420.110 1686.270 ;
        RECT 418.930 1683.490 420.110 1684.670 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -31.110 420.110 -29.930 ;
        RECT 418.930 -32.710 420.110 -31.530 ;
        RECT 598.930 3551.210 600.110 3552.390 ;
        RECT 598.930 3549.610 600.110 3550.790 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 598.930 3125.090 600.110 3126.270 ;
        RECT 598.930 3123.490 600.110 3124.670 ;
        RECT 598.930 2945.090 600.110 2946.270 ;
        RECT 598.930 2943.490 600.110 2944.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 598.930 2585.090 600.110 2586.270 ;
        RECT 598.930 2583.490 600.110 2584.670 ;
        RECT 598.930 2405.090 600.110 2406.270 ;
        RECT 598.930 2403.490 600.110 2404.670 ;
        RECT 598.930 2225.090 600.110 2226.270 ;
        RECT 598.930 2223.490 600.110 2224.670 ;
        RECT 598.930 2045.090 600.110 2046.270 ;
        RECT 598.930 2043.490 600.110 2044.670 ;
        RECT 598.930 1865.090 600.110 1866.270 ;
        RECT 598.930 1863.490 600.110 1864.670 ;
        RECT 598.930 1685.090 600.110 1686.270 ;
        RECT 598.930 1683.490 600.110 1684.670 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -31.110 600.110 -29.930 ;
        RECT 598.930 -32.710 600.110 -31.530 ;
        RECT 778.930 3551.210 780.110 3552.390 ;
        RECT 778.930 3549.610 780.110 3550.790 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 778.930 2585.090 780.110 2586.270 ;
        RECT 778.930 2583.490 780.110 2584.670 ;
        RECT 778.930 2405.090 780.110 2406.270 ;
        RECT 778.930 2403.490 780.110 2404.670 ;
        RECT 778.930 2225.090 780.110 2226.270 ;
        RECT 778.930 2223.490 780.110 2224.670 ;
        RECT 778.930 2045.090 780.110 2046.270 ;
        RECT 778.930 2043.490 780.110 2044.670 ;
        RECT 778.930 1865.090 780.110 1866.270 ;
        RECT 778.930 1863.490 780.110 1864.670 ;
        RECT 778.930 1685.090 780.110 1686.270 ;
        RECT 778.930 1683.490 780.110 1684.670 ;
        RECT 778.930 1505.090 780.110 1506.270 ;
        RECT 778.930 1503.490 780.110 1504.670 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 778.930 965.090 780.110 966.270 ;
        RECT 778.930 963.490 780.110 964.670 ;
        RECT 778.930 785.090 780.110 786.270 ;
        RECT 778.930 783.490 780.110 784.670 ;
        RECT 778.930 605.090 780.110 606.270 ;
        RECT 778.930 603.490 780.110 604.670 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -31.110 780.110 -29.930 ;
        RECT 778.930 -32.710 780.110 -31.530 ;
        RECT 958.930 3551.210 960.110 3552.390 ;
        RECT 958.930 3549.610 960.110 3550.790 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 958.930 3125.090 960.110 3126.270 ;
        RECT 958.930 3123.490 960.110 3124.670 ;
        RECT 958.930 2945.090 960.110 2946.270 ;
        RECT 958.930 2943.490 960.110 2944.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 958.930 2585.090 960.110 2586.270 ;
        RECT 958.930 2583.490 960.110 2584.670 ;
        RECT 958.930 2405.090 960.110 2406.270 ;
        RECT 958.930 2403.490 960.110 2404.670 ;
        RECT 958.930 2225.090 960.110 2226.270 ;
        RECT 958.930 2223.490 960.110 2224.670 ;
        RECT 958.930 2045.090 960.110 2046.270 ;
        RECT 958.930 2043.490 960.110 2044.670 ;
        RECT 958.930 1865.090 960.110 1866.270 ;
        RECT 958.930 1863.490 960.110 1864.670 ;
        RECT 958.930 1685.090 960.110 1686.270 ;
        RECT 958.930 1683.490 960.110 1684.670 ;
        RECT 958.930 1505.090 960.110 1506.270 ;
        RECT 958.930 1503.490 960.110 1504.670 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 958.930 965.090 960.110 966.270 ;
        RECT 958.930 963.490 960.110 964.670 ;
        RECT 958.930 785.090 960.110 786.270 ;
        RECT 958.930 783.490 960.110 784.670 ;
        RECT 958.930 605.090 960.110 606.270 ;
        RECT 958.930 603.490 960.110 604.670 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -31.110 960.110 -29.930 ;
        RECT 958.930 -32.710 960.110 -31.530 ;
        RECT 1138.930 3551.210 1140.110 3552.390 ;
        RECT 1138.930 3549.610 1140.110 3550.790 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1138.930 3125.090 1140.110 3126.270 ;
        RECT 1138.930 3123.490 1140.110 3124.670 ;
        RECT 1138.930 2945.090 1140.110 2946.270 ;
        RECT 1138.930 2943.490 1140.110 2944.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1138.930 2585.090 1140.110 2586.270 ;
        RECT 1138.930 2583.490 1140.110 2584.670 ;
        RECT 1138.930 2405.090 1140.110 2406.270 ;
        RECT 1138.930 2403.490 1140.110 2404.670 ;
        RECT 1138.930 2225.090 1140.110 2226.270 ;
        RECT 1138.930 2223.490 1140.110 2224.670 ;
        RECT 1138.930 2045.090 1140.110 2046.270 ;
        RECT 1138.930 2043.490 1140.110 2044.670 ;
        RECT 1138.930 1865.090 1140.110 1866.270 ;
        RECT 1138.930 1863.490 1140.110 1864.670 ;
        RECT 1138.930 1685.090 1140.110 1686.270 ;
        RECT 1138.930 1683.490 1140.110 1684.670 ;
        RECT 1138.930 1505.090 1140.110 1506.270 ;
        RECT 1138.930 1503.490 1140.110 1504.670 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1138.930 965.090 1140.110 966.270 ;
        RECT 1138.930 963.490 1140.110 964.670 ;
        RECT 1138.930 785.090 1140.110 786.270 ;
        RECT 1138.930 783.490 1140.110 784.670 ;
        RECT 1138.930 605.090 1140.110 606.270 ;
        RECT 1138.930 603.490 1140.110 604.670 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -31.110 1140.110 -29.930 ;
        RECT 1138.930 -32.710 1140.110 -31.530 ;
        RECT 1318.930 3551.210 1320.110 3552.390 ;
        RECT 1318.930 3549.610 1320.110 3550.790 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1318.930 3125.090 1320.110 3126.270 ;
        RECT 1318.930 3123.490 1320.110 3124.670 ;
        RECT 1318.930 2945.090 1320.110 2946.270 ;
        RECT 1318.930 2943.490 1320.110 2944.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1318.930 2585.090 1320.110 2586.270 ;
        RECT 1318.930 2583.490 1320.110 2584.670 ;
        RECT 1318.930 2405.090 1320.110 2406.270 ;
        RECT 1318.930 2403.490 1320.110 2404.670 ;
        RECT 1318.930 2225.090 1320.110 2226.270 ;
        RECT 1318.930 2223.490 1320.110 2224.670 ;
        RECT 1318.930 2045.090 1320.110 2046.270 ;
        RECT 1318.930 2043.490 1320.110 2044.670 ;
        RECT 1318.930 1865.090 1320.110 1866.270 ;
        RECT 1318.930 1863.490 1320.110 1864.670 ;
        RECT 1318.930 1685.090 1320.110 1686.270 ;
        RECT 1318.930 1683.490 1320.110 1684.670 ;
        RECT 1318.930 1505.090 1320.110 1506.270 ;
        RECT 1318.930 1503.490 1320.110 1504.670 ;
        RECT 1318.930 1325.090 1320.110 1326.270 ;
        RECT 1318.930 1323.490 1320.110 1324.670 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1318.930 965.090 1320.110 966.270 ;
        RECT 1318.930 963.490 1320.110 964.670 ;
        RECT 1318.930 785.090 1320.110 786.270 ;
        RECT 1318.930 783.490 1320.110 784.670 ;
        RECT 1318.930 605.090 1320.110 606.270 ;
        RECT 1318.930 603.490 1320.110 604.670 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -31.110 1320.110 -29.930 ;
        RECT 1318.930 -32.710 1320.110 -31.530 ;
        RECT 1498.930 3551.210 1500.110 3552.390 ;
        RECT 1498.930 3549.610 1500.110 3550.790 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 1498.930 2765.090 1500.110 2766.270 ;
        RECT 1498.930 2763.490 1500.110 2764.670 ;
        RECT 1498.930 2585.090 1500.110 2586.270 ;
        RECT 1498.930 2583.490 1500.110 2584.670 ;
        RECT 1498.930 2405.090 1500.110 2406.270 ;
        RECT 1498.930 2403.490 1500.110 2404.670 ;
        RECT 1498.930 2225.090 1500.110 2226.270 ;
        RECT 1498.930 2223.490 1500.110 2224.670 ;
        RECT 1498.930 2045.090 1500.110 2046.270 ;
        RECT 1498.930 2043.490 1500.110 2044.670 ;
        RECT 1498.930 1865.090 1500.110 1866.270 ;
        RECT 1498.930 1863.490 1500.110 1864.670 ;
        RECT 1498.930 1685.090 1500.110 1686.270 ;
        RECT 1498.930 1683.490 1500.110 1684.670 ;
        RECT 1498.930 1505.090 1500.110 1506.270 ;
        RECT 1498.930 1503.490 1500.110 1504.670 ;
        RECT 1498.930 1325.090 1500.110 1326.270 ;
        RECT 1498.930 1323.490 1500.110 1324.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1498.930 965.090 1500.110 966.270 ;
        RECT 1498.930 963.490 1500.110 964.670 ;
        RECT 1498.930 785.090 1500.110 786.270 ;
        RECT 1498.930 783.490 1500.110 784.670 ;
        RECT 1498.930 605.090 1500.110 606.270 ;
        RECT 1498.930 603.490 1500.110 604.670 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -31.110 1500.110 -29.930 ;
        RECT 1498.930 -32.710 1500.110 -31.530 ;
        RECT 1678.930 3551.210 1680.110 3552.390 ;
        RECT 1678.930 3549.610 1680.110 3550.790 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1678.930 2945.090 1680.110 2946.270 ;
        RECT 1678.930 2943.490 1680.110 2944.670 ;
        RECT 1678.930 2765.090 1680.110 2766.270 ;
        RECT 1678.930 2763.490 1680.110 2764.670 ;
        RECT 1678.930 2585.090 1680.110 2586.270 ;
        RECT 1678.930 2583.490 1680.110 2584.670 ;
        RECT 1678.930 2405.090 1680.110 2406.270 ;
        RECT 1678.930 2403.490 1680.110 2404.670 ;
        RECT 1678.930 2225.090 1680.110 2226.270 ;
        RECT 1678.930 2223.490 1680.110 2224.670 ;
        RECT 1678.930 2045.090 1680.110 2046.270 ;
        RECT 1678.930 2043.490 1680.110 2044.670 ;
        RECT 1678.930 1865.090 1680.110 1866.270 ;
        RECT 1678.930 1863.490 1680.110 1864.670 ;
        RECT 1678.930 1685.090 1680.110 1686.270 ;
        RECT 1678.930 1683.490 1680.110 1684.670 ;
        RECT 1678.930 1505.090 1680.110 1506.270 ;
        RECT 1678.930 1503.490 1680.110 1504.670 ;
        RECT 1678.930 1325.090 1680.110 1326.270 ;
        RECT 1678.930 1323.490 1680.110 1324.670 ;
        RECT 1678.930 1145.090 1680.110 1146.270 ;
        RECT 1678.930 1143.490 1680.110 1144.670 ;
        RECT 1678.930 965.090 1680.110 966.270 ;
        RECT 1678.930 963.490 1680.110 964.670 ;
        RECT 1678.930 785.090 1680.110 786.270 ;
        RECT 1678.930 783.490 1680.110 784.670 ;
        RECT 1678.930 605.090 1680.110 606.270 ;
        RECT 1678.930 603.490 1680.110 604.670 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -31.110 1680.110 -29.930 ;
        RECT 1678.930 -32.710 1680.110 -31.530 ;
        RECT 1858.930 3551.210 1860.110 3552.390 ;
        RECT 1858.930 3549.610 1860.110 3550.790 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 1858.930 2945.090 1860.110 2946.270 ;
        RECT 1858.930 2943.490 1860.110 2944.670 ;
        RECT 1858.930 2765.090 1860.110 2766.270 ;
        RECT 1858.930 2763.490 1860.110 2764.670 ;
        RECT 1858.930 2585.090 1860.110 2586.270 ;
        RECT 1858.930 2583.490 1860.110 2584.670 ;
        RECT 1858.930 2405.090 1860.110 2406.270 ;
        RECT 1858.930 2403.490 1860.110 2404.670 ;
        RECT 1858.930 2225.090 1860.110 2226.270 ;
        RECT 1858.930 2223.490 1860.110 2224.670 ;
        RECT 1858.930 2045.090 1860.110 2046.270 ;
        RECT 1858.930 2043.490 1860.110 2044.670 ;
        RECT 1858.930 1865.090 1860.110 1866.270 ;
        RECT 1858.930 1863.490 1860.110 1864.670 ;
        RECT 1858.930 1685.090 1860.110 1686.270 ;
        RECT 1858.930 1683.490 1860.110 1684.670 ;
        RECT 1858.930 1505.090 1860.110 1506.270 ;
        RECT 1858.930 1503.490 1860.110 1504.670 ;
        RECT 1858.930 1325.090 1860.110 1326.270 ;
        RECT 1858.930 1323.490 1860.110 1324.670 ;
        RECT 1858.930 1145.090 1860.110 1146.270 ;
        RECT 1858.930 1143.490 1860.110 1144.670 ;
        RECT 1858.930 965.090 1860.110 966.270 ;
        RECT 1858.930 963.490 1860.110 964.670 ;
        RECT 1858.930 785.090 1860.110 786.270 ;
        RECT 1858.930 783.490 1860.110 784.670 ;
        RECT 1858.930 605.090 1860.110 606.270 ;
        RECT 1858.930 603.490 1860.110 604.670 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -31.110 1860.110 -29.930 ;
        RECT 1858.930 -32.710 1860.110 -31.530 ;
        RECT 2038.930 3551.210 2040.110 3552.390 ;
        RECT 2038.930 3549.610 2040.110 3550.790 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 2038.930 2405.090 2040.110 2406.270 ;
        RECT 2038.930 2403.490 2040.110 2404.670 ;
        RECT 2038.930 2225.090 2040.110 2226.270 ;
        RECT 2038.930 2223.490 2040.110 2224.670 ;
        RECT 2038.930 2045.090 2040.110 2046.270 ;
        RECT 2038.930 2043.490 2040.110 2044.670 ;
        RECT 2038.930 1865.090 2040.110 1866.270 ;
        RECT 2038.930 1863.490 2040.110 1864.670 ;
        RECT 2038.930 1685.090 2040.110 1686.270 ;
        RECT 2038.930 1683.490 2040.110 1684.670 ;
        RECT 2038.930 1505.090 2040.110 1506.270 ;
        RECT 2038.930 1503.490 2040.110 1504.670 ;
        RECT 2038.930 1325.090 2040.110 1326.270 ;
        RECT 2038.930 1323.490 2040.110 1324.670 ;
        RECT 2038.930 1145.090 2040.110 1146.270 ;
        RECT 2038.930 1143.490 2040.110 1144.670 ;
        RECT 2038.930 965.090 2040.110 966.270 ;
        RECT 2038.930 963.490 2040.110 964.670 ;
        RECT 2038.930 785.090 2040.110 786.270 ;
        RECT 2038.930 783.490 2040.110 784.670 ;
        RECT 2038.930 605.090 2040.110 606.270 ;
        RECT 2038.930 603.490 2040.110 604.670 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -31.110 2040.110 -29.930 ;
        RECT 2038.930 -32.710 2040.110 -31.530 ;
        RECT 2218.930 3551.210 2220.110 3552.390 ;
        RECT 2218.930 3549.610 2220.110 3550.790 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2218.930 2945.090 2220.110 2946.270 ;
        RECT 2218.930 2943.490 2220.110 2944.670 ;
        RECT 2218.930 2765.090 2220.110 2766.270 ;
        RECT 2218.930 2763.490 2220.110 2764.670 ;
        RECT 2218.930 2585.090 2220.110 2586.270 ;
        RECT 2218.930 2583.490 2220.110 2584.670 ;
        RECT 2218.930 2405.090 2220.110 2406.270 ;
        RECT 2218.930 2403.490 2220.110 2404.670 ;
        RECT 2218.930 2225.090 2220.110 2226.270 ;
        RECT 2218.930 2223.490 2220.110 2224.670 ;
        RECT 2218.930 2045.090 2220.110 2046.270 ;
        RECT 2218.930 2043.490 2220.110 2044.670 ;
        RECT 2218.930 1865.090 2220.110 1866.270 ;
        RECT 2218.930 1863.490 2220.110 1864.670 ;
        RECT 2218.930 1685.090 2220.110 1686.270 ;
        RECT 2218.930 1683.490 2220.110 1684.670 ;
        RECT 2218.930 1505.090 2220.110 1506.270 ;
        RECT 2218.930 1503.490 2220.110 1504.670 ;
        RECT 2218.930 1325.090 2220.110 1326.270 ;
        RECT 2218.930 1323.490 2220.110 1324.670 ;
        RECT 2218.930 1145.090 2220.110 1146.270 ;
        RECT 2218.930 1143.490 2220.110 1144.670 ;
        RECT 2218.930 965.090 2220.110 966.270 ;
        RECT 2218.930 963.490 2220.110 964.670 ;
        RECT 2218.930 785.090 2220.110 786.270 ;
        RECT 2218.930 783.490 2220.110 784.670 ;
        RECT 2218.930 605.090 2220.110 606.270 ;
        RECT 2218.930 603.490 2220.110 604.670 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -31.110 2220.110 -29.930 ;
        RECT 2218.930 -32.710 2220.110 -31.530 ;
        RECT 2398.930 3551.210 2400.110 3552.390 ;
        RECT 2398.930 3549.610 2400.110 3550.790 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2398.930 2945.090 2400.110 2946.270 ;
        RECT 2398.930 2943.490 2400.110 2944.670 ;
        RECT 2398.930 2765.090 2400.110 2766.270 ;
        RECT 2398.930 2763.490 2400.110 2764.670 ;
        RECT 2398.930 2585.090 2400.110 2586.270 ;
        RECT 2398.930 2583.490 2400.110 2584.670 ;
        RECT 2398.930 2405.090 2400.110 2406.270 ;
        RECT 2398.930 2403.490 2400.110 2404.670 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2398.930 2045.090 2400.110 2046.270 ;
        RECT 2398.930 2043.490 2400.110 2044.670 ;
        RECT 2398.930 1865.090 2400.110 1866.270 ;
        RECT 2398.930 1863.490 2400.110 1864.670 ;
        RECT 2398.930 1685.090 2400.110 1686.270 ;
        RECT 2398.930 1683.490 2400.110 1684.670 ;
        RECT 2398.930 1505.090 2400.110 1506.270 ;
        RECT 2398.930 1503.490 2400.110 1504.670 ;
        RECT 2398.930 1325.090 2400.110 1326.270 ;
        RECT 2398.930 1323.490 2400.110 1324.670 ;
        RECT 2398.930 1145.090 2400.110 1146.270 ;
        RECT 2398.930 1143.490 2400.110 1144.670 ;
        RECT 2398.930 965.090 2400.110 966.270 ;
        RECT 2398.930 963.490 2400.110 964.670 ;
        RECT 2398.930 785.090 2400.110 786.270 ;
        RECT 2398.930 783.490 2400.110 784.670 ;
        RECT 2398.930 605.090 2400.110 606.270 ;
        RECT 2398.930 603.490 2400.110 604.670 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -31.110 2400.110 -29.930 ;
        RECT 2398.930 -32.710 2400.110 -31.530 ;
        RECT 2578.930 3551.210 2580.110 3552.390 ;
        RECT 2578.930 3549.610 2580.110 3550.790 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -31.110 2580.110 -29.930 ;
        RECT 2578.930 -32.710 2580.110 -31.530 ;
        RECT 2758.930 3551.210 2760.110 3552.390 ;
        RECT 2758.930 3549.610 2760.110 3550.790 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -31.110 2760.110 -29.930 ;
        RECT 2758.930 -32.710 2760.110 -31.530 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT 2955.710 3485.090 2956.890 3486.270 ;
        RECT 2955.710 3483.490 2956.890 3484.670 ;
        RECT 2955.710 3305.090 2956.890 3306.270 ;
        RECT 2955.710 3303.490 2956.890 3304.670 ;
        RECT 2955.710 3125.090 2956.890 3126.270 ;
        RECT 2955.710 3123.490 2956.890 3124.670 ;
        RECT 2955.710 2945.090 2956.890 2946.270 ;
        RECT 2955.710 2943.490 2956.890 2944.670 ;
        RECT 2955.710 2765.090 2956.890 2766.270 ;
        RECT 2955.710 2763.490 2956.890 2764.670 ;
        RECT 2955.710 2585.090 2956.890 2586.270 ;
        RECT 2955.710 2583.490 2956.890 2584.670 ;
        RECT 2955.710 2405.090 2956.890 2406.270 ;
        RECT 2955.710 2403.490 2956.890 2404.670 ;
        RECT 2955.710 2225.090 2956.890 2226.270 ;
        RECT 2955.710 2223.490 2956.890 2224.670 ;
        RECT 2955.710 2045.090 2956.890 2046.270 ;
        RECT 2955.710 2043.490 2956.890 2044.670 ;
        RECT 2955.710 1865.090 2956.890 1866.270 ;
        RECT 2955.710 1863.490 2956.890 1864.670 ;
        RECT 2955.710 1685.090 2956.890 1686.270 ;
        RECT 2955.710 1683.490 2956.890 1684.670 ;
        RECT 2955.710 1505.090 2956.890 1506.270 ;
        RECT 2955.710 1503.490 2956.890 1504.670 ;
        RECT 2955.710 1325.090 2956.890 1326.270 ;
        RECT 2955.710 1323.490 2956.890 1324.670 ;
        RECT 2955.710 1145.090 2956.890 1146.270 ;
        RECT 2955.710 1143.490 2956.890 1144.670 ;
        RECT 2955.710 965.090 2956.890 966.270 ;
        RECT 2955.710 963.490 2956.890 964.670 ;
        RECT 2955.710 785.090 2956.890 786.270 ;
        RECT 2955.710 783.490 2956.890 784.670 ;
        RECT 2955.710 605.090 2956.890 606.270 ;
        RECT 2955.710 603.490 2956.890 604.670 ;
        RECT 2955.710 425.090 2956.890 426.270 ;
        RECT 2955.710 423.490 2956.890 424.670 ;
        RECT 2955.710 245.090 2956.890 246.270 ;
        RECT 2955.710 243.490 2956.890 244.670 ;
        RECT 2955.710 65.090 2956.890 66.270 ;
        RECT 2955.710 63.490 2956.890 64.670 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 58.020 3552.500 61.020 3552.510 ;
        RECT 238.020 3552.500 241.020 3552.510 ;
        RECT 418.020 3552.500 421.020 3552.510 ;
        RECT 598.020 3552.500 601.020 3552.510 ;
        RECT 778.020 3552.500 781.020 3552.510 ;
        RECT 958.020 3552.500 961.020 3552.510 ;
        RECT 1138.020 3552.500 1141.020 3552.510 ;
        RECT 1318.020 3552.500 1321.020 3552.510 ;
        RECT 1498.020 3552.500 1501.020 3552.510 ;
        RECT 1678.020 3552.500 1681.020 3552.510 ;
        RECT 1858.020 3552.500 1861.020 3552.510 ;
        RECT 2038.020 3552.500 2041.020 3552.510 ;
        RECT 2218.020 3552.500 2221.020 3552.510 ;
        RECT 2398.020 3552.500 2401.020 3552.510 ;
        RECT 2578.020 3552.500 2581.020 3552.510 ;
        RECT 2758.020 3552.500 2761.020 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 58.020 3549.490 61.020 3549.500 ;
        RECT 238.020 3549.490 241.020 3549.500 ;
        RECT 418.020 3549.490 421.020 3549.500 ;
        RECT 598.020 3549.490 601.020 3549.500 ;
        RECT 778.020 3549.490 781.020 3549.500 ;
        RECT 958.020 3549.490 961.020 3549.500 ;
        RECT 1138.020 3549.490 1141.020 3549.500 ;
        RECT 1318.020 3549.490 1321.020 3549.500 ;
        RECT 1498.020 3549.490 1501.020 3549.500 ;
        RECT 1678.020 3549.490 1681.020 3549.500 ;
        RECT 1858.020 3549.490 1861.020 3549.500 ;
        RECT 2038.020 3549.490 2041.020 3549.500 ;
        RECT 2218.020 3549.490 2221.020 3549.500 ;
        RECT 2398.020 3549.490 2401.020 3549.500 ;
        RECT 2578.020 3549.490 2581.020 3549.500 ;
        RECT 2758.020 3549.490 2761.020 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -38.180 3486.380 -35.180 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.800 3486.380 2957.800 3486.390 ;
        RECT -42.880 3483.380 2962.500 3486.380 ;
        RECT -38.180 3483.370 -35.180 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.800 3483.370 2957.800 3483.380 ;
        RECT -38.180 3306.380 -35.180 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.800 3306.380 2957.800 3306.390 ;
        RECT -42.880 3303.380 2962.500 3306.380 ;
        RECT -38.180 3303.370 -35.180 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.800 3303.370 2957.800 3303.380 ;
        RECT -38.180 3126.380 -35.180 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 418.020 3126.380 421.020 3126.390 ;
        RECT 598.020 3126.380 601.020 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 958.020 3126.380 961.020 3126.390 ;
        RECT 1138.020 3126.380 1141.020 3126.390 ;
        RECT 1318.020 3126.380 1321.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.800 3126.380 2957.800 3126.390 ;
        RECT -42.880 3123.380 2962.500 3126.380 ;
        RECT -38.180 3123.370 -35.180 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 418.020 3123.370 421.020 3123.380 ;
        RECT 598.020 3123.370 601.020 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 958.020 3123.370 961.020 3123.380 ;
        RECT 1138.020 3123.370 1141.020 3123.380 ;
        RECT 1318.020 3123.370 1321.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.800 3123.370 2957.800 3123.380 ;
        RECT -38.180 2946.380 -35.180 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 418.020 2946.380 421.020 2946.390 ;
        RECT 598.020 2946.380 601.020 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 958.020 2946.380 961.020 2946.390 ;
        RECT 1138.020 2946.380 1141.020 2946.390 ;
        RECT 1318.020 2946.380 1321.020 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1678.020 2946.380 1681.020 2946.390 ;
        RECT 1858.020 2946.380 1861.020 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2218.020 2946.380 2221.020 2946.390 ;
        RECT 2398.020 2946.380 2401.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.800 2946.380 2957.800 2946.390 ;
        RECT -42.880 2943.380 2962.500 2946.380 ;
        RECT -38.180 2943.370 -35.180 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 418.020 2943.370 421.020 2943.380 ;
        RECT 598.020 2943.370 601.020 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 958.020 2943.370 961.020 2943.380 ;
        RECT 1138.020 2943.370 1141.020 2943.380 ;
        RECT 1318.020 2943.370 1321.020 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1678.020 2943.370 1681.020 2943.380 ;
        RECT 1858.020 2943.370 1861.020 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2218.020 2943.370 2221.020 2943.380 ;
        RECT 2398.020 2943.370 2401.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.800 2943.370 2957.800 2943.380 ;
        RECT -38.180 2766.380 -35.180 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 1498.020 2766.380 1501.020 2766.390 ;
        RECT 1678.020 2766.380 1681.020 2766.390 ;
        RECT 1858.020 2766.380 1861.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2218.020 2766.380 2221.020 2766.390 ;
        RECT 2398.020 2766.380 2401.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.800 2766.380 2957.800 2766.390 ;
        RECT -42.880 2763.380 2962.500 2766.380 ;
        RECT -38.180 2763.370 -35.180 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 1498.020 2763.370 1501.020 2763.380 ;
        RECT 1678.020 2763.370 1681.020 2763.380 ;
        RECT 1858.020 2763.370 1861.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2218.020 2763.370 2221.020 2763.380 ;
        RECT 2398.020 2763.370 2401.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.800 2763.370 2957.800 2763.380 ;
        RECT -38.180 2586.380 -35.180 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 418.020 2586.380 421.020 2586.390 ;
        RECT 598.020 2586.380 601.020 2586.390 ;
        RECT 778.020 2586.380 781.020 2586.390 ;
        RECT 958.020 2586.380 961.020 2586.390 ;
        RECT 1138.020 2586.380 1141.020 2586.390 ;
        RECT 1318.020 2586.380 1321.020 2586.390 ;
        RECT 1498.020 2586.380 1501.020 2586.390 ;
        RECT 1678.020 2586.380 1681.020 2586.390 ;
        RECT 1858.020 2586.380 1861.020 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2218.020 2586.380 2221.020 2586.390 ;
        RECT 2398.020 2586.380 2401.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.800 2586.380 2957.800 2586.390 ;
        RECT -42.880 2583.380 2962.500 2586.380 ;
        RECT -38.180 2583.370 -35.180 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 418.020 2583.370 421.020 2583.380 ;
        RECT 598.020 2583.370 601.020 2583.380 ;
        RECT 778.020 2583.370 781.020 2583.380 ;
        RECT 958.020 2583.370 961.020 2583.380 ;
        RECT 1138.020 2583.370 1141.020 2583.380 ;
        RECT 1318.020 2583.370 1321.020 2583.380 ;
        RECT 1498.020 2583.370 1501.020 2583.380 ;
        RECT 1678.020 2583.370 1681.020 2583.380 ;
        RECT 1858.020 2583.370 1861.020 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2218.020 2583.370 2221.020 2583.380 ;
        RECT 2398.020 2583.370 2401.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.800 2583.370 2957.800 2583.380 ;
        RECT -38.180 2406.380 -35.180 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 418.020 2406.380 421.020 2406.390 ;
        RECT 598.020 2406.380 601.020 2406.390 ;
        RECT 778.020 2406.380 781.020 2406.390 ;
        RECT 958.020 2406.380 961.020 2406.390 ;
        RECT 1138.020 2406.380 1141.020 2406.390 ;
        RECT 1318.020 2406.380 1321.020 2406.390 ;
        RECT 1498.020 2406.380 1501.020 2406.390 ;
        RECT 1678.020 2406.380 1681.020 2406.390 ;
        RECT 1858.020 2406.380 1861.020 2406.390 ;
        RECT 2038.020 2406.380 2041.020 2406.390 ;
        RECT 2218.020 2406.380 2221.020 2406.390 ;
        RECT 2398.020 2406.380 2401.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.800 2406.380 2957.800 2406.390 ;
        RECT -42.880 2403.380 2962.500 2406.380 ;
        RECT -38.180 2403.370 -35.180 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 418.020 2403.370 421.020 2403.380 ;
        RECT 598.020 2403.370 601.020 2403.380 ;
        RECT 778.020 2403.370 781.020 2403.380 ;
        RECT 958.020 2403.370 961.020 2403.380 ;
        RECT 1138.020 2403.370 1141.020 2403.380 ;
        RECT 1318.020 2403.370 1321.020 2403.380 ;
        RECT 1498.020 2403.370 1501.020 2403.380 ;
        RECT 1678.020 2403.370 1681.020 2403.380 ;
        RECT 1858.020 2403.370 1861.020 2403.380 ;
        RECT 2038.020 2403.370 2041.020 2403.380 ;
        RECT 2218.020 2403.370 2221.020 2403.380 ;
        RECT 2398.020 2403.370 2401.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.800 2403.370 2957.800 2403.380 ;
        RECT -38.180 2226.380 -35.180 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 418.020 2226.380 421.020 2226.390 ;
        RECT 598.020 2226.380 601.020 2226.390 ;
        RECT 778.020 2226.380 781.020 2226.390 ;
        RECT 958.020 2226.380 961.020 2226.390 ;
        RECT 1138.020 2226.380 1141.020 2226.390 ;
        RECT 1318.020 2226.380 1321.020 2226.390 ;
        RECT 1498.020 2226.380 1501.020 2226.390 ;
        RECT 1678.020 2226.380 1681.020 2226.390 ;
        RECT 1858.020 2226.380 1861.020 2226.390 ;
        RECT 2038.020 2226.380 2041.020 2226.390 ;
        RECT 2218.020 2226.380 2221.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.800 2226.380 2957.800 2226.390 ;
        RECT -42.880 2223.380 2962.500 2226.380 ;
        RECT -38.180 2223.370 -35.180 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 418.020 2223.370 421.020 2223.380 ;
        RECT 598.020 2223.370 601.020 2223.380 ;
        RECT 778.020 2223.370 781.020 2223.380 ;
        RECT 958.020 2223.370 961.020 2223.380 ;
        RECT 1138.020 2223.370 1141.020 2223.380 ;
        RECT 1318.020 2223.370 1321.020 2223.380 ;
        RECT 1498.020 2223.370 1501.020 2223.380 ;
        RECT 1678.020 2223.370 1681.020 2223.380 ;
        RECT 1858.020 2223.370 1861.020 2223.380 ;
        RECT 2038.020 2223.370 2041.020 2223.380 ;
        RECT 2218.020 2223.370 2221.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.800 2223.370 2957.800 2223.380 ;
        RECT -38.180 2046.380 -35.180 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 418.020 2046.380 421.020 2046.390 ;
        RECT 598.020 2046.380 601.020 2046.390 ;
        RECT 778.020 2046.380 781.020 2046.390 ;
        RECT 958.020 2046.380 961.020 2046.390 ;
        RECT 1138.020 2046.380 1141.020 2046.390 ;
        RECT 1318.020 2046.380 1321.020 2046.390 ;
        RECT 1498.020 2046.380 1501.020 2046.390 ;
        RECT 1678.020 2046.380 1681.020 2046.390 ;
        RECT 1858.020 2046.380 1861.020 2046.390 ;
        RECT 2038.020 2046.380 2041.020 2046.390 ;
        RECT 2218.020 2046.380 2221.020 2046.390 ;
        RECT 2398.020 2046.380 2401.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.800 2046.380 2957.800 2046.390 ;
        RECT -42.880 2043.380 2962.500 2046.380 ;
        RECT -38.180 2043.370 -35.180 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 418.020 2043.370 421.020 2043.380 ;
        RECT 598.020 2043.370 601.020 2043.380 ;
        RECT 778.020 2043.370 781.020 2043.380 ;
        RECT 958.020 2043.370 961.020 2043.380 ;
        RECT 1138.020 2043.370 1141.020 2043.380 ;
        RECT 1318.020 2043.370 1321.020 2043.380 ;
        RECT 1498.020 2043.370 1501.020 2043.380 ;
        RECT 1678.020 2043.370 1681.020 2043.380 ;
        RECT 1858.020 2043.370 1861.020 2043.380 ;
        RECT 2038.020 2043.370 2041.020 2043.380 ;
        RECT 2218.020 2043.370 2221.020 2043.380 ;
        RECT 2398.020 2043.370 2401.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.800 2043.370 2957.800 2043.380 ;
        RECT -38.180 1866.380 -35.180 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 418.020 1866.380 421.020 1866.390 ;
        RECT 598.020 1866.380 601.020 1866.390 ;
        RECT 778.020 1866.380 781.020 1866.390 ;
        RECT 958.020 1866.380 961.020 1866.390 ;
        RECT 1138.020 1866.380 1141.020 1866.390 ;
        RECT 1318.020 1866.380 1321.020 1866.390 ;
        RECT 1498.020 1866.380 1501.020 1866.390 ;
        RECT 1678.020 1866.380 1681.020 1866.390 ;
        RECT 1858.020 1866.380 1861.020 1866.390 ;
        RECT 2038.020 1866.380 2041.020 1866.390 ;
        RECT 2218.020 1866.380 2221.020 1866.390 ;
        RECT 2398.020 1866.380 2401.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.800 1866.380 2957.800 1866.390 ;
        RECT -42.880 1863.380 2962.500 1866.380 ;
        RECT -38.180 1863.370 -35.180 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 418.020 1863.370 421.020 1863.380 ;
        RECT 598.020 1863.370 601.020 1863.380 ;
        RECT 778.020 1863.370 781.020 1863.380 ;
        RECT 958.020 1863.370 961.020 1863.380 ;
        RECT 1138.020 1863.370 1141.020 1863.380 ;
        RECT 1318.020 1863.370 1321.020 1863.380 ;
        RECT 1498.020 1863.370 1501.020 1863.380 ;
        RECT 1678.020 1863.370 1681.020 1863.380 ;
        RECT 1858.020 1863.370 1861.020 1863.380 ;
        RECT 2038.020 1863.370 2041.020 1863.380 ;
        RECT 2218.020 1863.370 2221.020 1863.380 ;
        RECT 2398.020 1863.370 2401.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.800 1863.370 2957.800 1863.380 ;
        RECT -38.180 1686.380 -35.180 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 418.020 1686.380 421.020 1686.390 ;
        RECT 598.020 1686.380 601.020 1686.390 ;
        RECT 778.020 1686.380 781.020 1686.390 ;
        RECT 958.020 1686.380 961.020 1686.390 ;
        RECT 1138.020 1686.380 1141.020 1686.390 ;
        RECT 1318.020 1686.380 1321.020 1686.390 ;
        RECT 1498.020 1686.380 1501.020 1686.390 ;
        RECT 1678.020 1686.380 1681.020 1686.390 ;
        RECT 1858.020 1686.380 1861.020 1686.390 ;
        RECT 2038.020 1686.380 2041.020 1686.390 ;
        RECT 2218.020 1686.380 2221.020 1686.390 ;
        RECT 2398.020 1686.380 2401.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.800 1686.380 2957.800 1686.390 ;
        RECT -42.880 1683.380 2962.500 1686.380 ;
        RECT -38.180 1683.370 -35.180 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 418.020 1683.370 421.020 1683.380 ;
        RECT 598.020 1683.370 601.020 1683.380 ;
        RECT 778.020 1683.370 781.020 1683.380 ;
        RECT 958.020 1683.370 961.020 1683.380 ;
        RECT 1138.020 1683.370 1141.020 1683.380 ;
        RECT 1318.020 1683.370 1321.020 1683.380 ;
        RECT 1498.020 1683.370 1501.020 1683.380 ;
        RECT 1678.020 1683.370 1681.020 1683.380 ;
        RECT 1858.020 1683.370 1861.020 1683.380 ;
        RECT 2038.020 1683.370 2041.020 1683.380 ;
        RECT 2218.020 1683.370 2221.020 1683.380 ;
        RECT 2398.020 1683.370 2401.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.800 1683.370 2957.800 1683.380 ;
        RECT -38.180 1506.380 -35.180 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 778.020 1506.380 781.020 1506.390 ;
        RECT 958.020 1506.380 961.020 1506.390 ;
        RECT 1138.020 1506.380 1141.020 1506.390 ;
        RECT 1318.020 1506.380 1321.020 1506.390 ;
        RECT 1498.020 1506.380 1501.020 1506.390 ;
        RECT 1678.020 1506.380 1681.020 1506.390 ;
        RECT 1858.020 1506.380 1861.020 1506.390 ;
        RECT 2038.020 1506.380 2041.020 1506.390 ;
        RECT 2218.020 1506.380 2221.020 1506.390 ;
        RECT 2398.020 1506.380 2401.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.800 1506.380 2957.800 1506.390 ;
        RECT -42.880 1503.380 2962.500 1506.380 ;
        RECT -38.180 1503.370 -35.180 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 778.020 1503.370 781.020 1503.380 ;
        RECT 958.020 1503.370 961.020 1503.380 ;
        RECT 1138.020 1503.370 1141.020 1503.380 ;
        RECT 1318.020 1503.370 1321.020 1503.380 ;
        RECT 1498.020 1503.370 1501.020 1503.380 ;
        RECT 1678.020 1503.370 1681.020 1503.380 ;
        RECT 1858.020 1503.370 1861.020 1503.380 ;
        RECT 2038.020 1503.370 2041.020 1503.380 ;
        RECT 2218.020 1503.370 2221.020 1503.380 ;
        RECT 2398.020 1503.370 2401.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.800 1503.370 2957.800 1503.380 ;
        RECT -38.180 1326.380 -35.180 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 1318.020 1326.380 1321.020 1326.390 ;
        RECT 1498.020 1326.380 1501.020 1326.390 ;
        RECT 1678.020 1326.380 1681.020 1326.390 ;
        RECT 1858.020 1326.380 1861.020 1326.390 ;
        RECT 2038.020 1326.380 2041.020 1326.390 ;
        RECT 2218.020 1326.380 2221.020 1326.390 ;
        RECT 2398.020 1326.380 2401.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.800 1326.380 2957.800 1326.390 ;
        RECT -42.880 1323.380 2962.500 1326.380 ;
        RECT -38.180 1323.370 -35.180 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 1318.020 1323.370 1321.020 1323.380 ;
        RECT 1498.020 1323.370 1501.020 1323.380 ;
        RECT 1678.020 1323.370 1681.020 1323.380 ;
        RECT 1858.020 1323.370 1861.020 1323.380 ;
        RECT 2038.020 1323.370 2041.020 1323.380 ;
        RECT 2218.020 1323.370 2221.020 1323.380 ;
        RECT 2398.020 1323.370 2401.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.800 1323.370 2957.800 1323.380 ;
        RECT -38.180 1146.380 -35.180 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1678.020 1146.380 1681.020 1146.390 ;
        RECT 1858.020 1146.380 1861.020 1146.390 ;
        RECT 2038.020 1146.380 2041.020 1146.390 ;
        RECT 2218.020 1146.380 2221.020 1146.390 ;
        RECT 2398.020 1146.380 2401.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.800 1146.380 2957.800 1146.390 ;
        RECT -42.880 1143.380 2962.500 1146.380 ;
        RECT -38.180 1143.370 -35.180 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1678.020 1143.370 1681.020 1143.380 ;
        RECT 1858.020 1143.370 1861.020 1143.380 ;
        RECT 2038.020 1143.370 2041.020 1143.380 ;
        RECT 2218.020 1143.370 2221.020 1143.380 ;
        RECT 2398.020 1143.370 2401.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.800 1143.370 2957.800 1143.380 ;
        RECT -38.180 966.380 -35.180 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 778.020 966.380 781.020 966.390 ;
        RECT 958.020 966.380 961.020 966.390 ;
        RECT 1138.020 966.380 1141.020 966.390 ;
        RECT 1318.020 966.380 1321.020 966.390 ;
        RECT 1498.020 966.380 1501.020 966.390 ;
        RECT 1678.020 966.380 1681.020 966.390 ;
        RECT 1858.020 966.380 1861.020 966.390 ;
        RECT 2038.020 966.380 2041.020 966.390 ;
        RECT 2218.020 966.380 2221.020 966.390 ;
        RECT 2398.020 966.380 2401.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.800 966.380 2957.800 966.390 ;
        RECT -42.880 963.380 2962.500 966.380 ;
        RECT -38.180 963.370 -35.180 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 778.020 963.370 781.020 963.380 ;
        RECT 958.020 963.370 961.020 963.380 ;
        RECT 1138.020 963.370 1141.020 963.380 ;
        RECT 1318.020 963.370 1321.020 963.380 ;
        RECT 1498.020 963.370 1501.020 963.380 ;
        RECT 1678.020 963.370 1681.020 963.380 ;
        RECT 1858.020 963.370 1861.020 963.380 ;
        RECT 2038.020 963.370 2041.020 963.380 ;
        RECT 2218.020 963.370 2221.020 963.380 ;
        RECT 2398.020 963.370 2401.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.800 963.370 2957.800 963.380 ;
        RECT -38.180 786.380 -35.180 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 778.020 786.380 781.020 786.390 ;
        RECT 958.020 786.380 961.020 786.390 ;
        RECT 1138.020 786.380 1141.020 786.390 ;
        RECT 1318.020 786.380 1321.020 786.390 ;
        RECT 1498.020 786.380 1501.020 786.390 ;
        RECT 1678.020 786.380 1681.020 786.390 ;
        RECT 1858.020 786.380 1861.020 786.390 ;
        RECT 2038.020 786.380 2041.020 786.390 ;
        RECT 2218.020 786.380 2221.020 786.390 ;
        RECT 2398.020 786.380 2401.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.800 786.380 2957.800 786.390 ;
        RECT -42.880 783.380 2962.500 786.380 ;
        RECT -38.180 783.370 -35.180 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 778.020 783.370 781.020 783.380 ;
        RECT 958.020 783.370 961.020 783.380 ;
        RECT 1138.020 783.370 1141.020 783.380 ;
        RECT 1318.020 783.370 1321.020 783.380 ;
        RECT 1498.020 783.370 1501.020 783.380 ;
        RECT 1678.020 783.370 1681.020 783.380 ;
        RECT 1858.020 783.370 1861.020 783.380 ;
        RECT 2038.020 783.370 2041.020 783.380 ;
        RECT 2218.020 783.370 2221.020 783.380 ;
        RECT 2398.020 783.370 2401.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.800 783.370 2957.800 783.380 ;
        RECT -38.180 606.380 -35.180 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 778.020 606.380 781.020 606.390 ;
        RECT 958.020 606.380 961.020 606.390 ;
        RECT 1138.020 606.380 1141.020 606.390 ;
        RECT 1318.020 606.380 1321.020 606.390 ;
        RECT 1498.020 606.380 1501.020 606.390 ;
        RECT 1678.020 606.380 1681.020 606.390 ;
        RECT 1858.020 606.380 1861.020 606.390 ;
        RECT 2038.020 606.380 2041.020 606.390 ;
        RECT 2218.020 606.380 2221.020 606.390 ;
        RECT 2398.020 606.380 2401.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.800 606.380 2957.800 606.390 ;
        RECT -42.880 603.380 2962.500 606.380 ;
        RECT -38.180 603.370 -35.180 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 778.020 603.370 781.020 603.380 ;
        RECT 958.020 603.370 961.020 603.380 ;
        RECT 1138.020 603.370 1141.020 603.380 ;
        RECT 1318.020 603.370 1321.020 603.380 ;
        RECT 1498.020 603.370 1501.020 603.380 ;
        RECT 1678.020 603.370 1681.020 603.380 ;
        RECT 1858.020 603.370 1861.020 603.380 ;
        RECT 2038.020 603.370 2041.020 603.380 ;
        RECT 2218.020 603.370 2221.020 603.380 ;
        RECT 2398.020 603.370 2401.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.800 603.370 2957.800 603.380 ;
        RECT -38.180 426.380 -35.180 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.800 426.380 2957.800 426.390 ;
        RECT -42.880 423.380 2962.500 426.380 ;
        RECT -38.180 423.370 -35.180 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.800 423.370 2957.800 423.380 ;
        RECT -38.180 246.380 -35.180 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.800 246.380 2957.800 246.390 ;
        RECT -42.880 243.380 2962.500 246.380 ;
        RECT -38.180 243.370 -35.180 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.800 243.370 2957.800 243.380 ;
        RECT -38.180 66.380 -35.180 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.800 66.380 2957.800 66.390 ;
        RECT -42.880 63.380 2962.500 66.380 ;
        RECT -38.180 63.370 -35.180 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.800 63.370 2957.800 63.380 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 58.020 -29.820 61.020 -29.810 ;
        RECT 238.020 -29.820 241.020 -29.810 ;
        RECT 418.020 -29.820 421.020 -29.810 ;
        RECT 598.020 -29.820 601.020 -29.810 ;
        RECT 778.020 -29.820 781.020 -29.810 ;
        RECT 958.020 -29.820 961.020 -29.810 ;
        RECT 1138.020 -29.820 1141.020 -29.810 ;
        RECT 1318.020 -29.820 1321.020 -29.810 ;
        RECT 1498.020 -29.820 1501.020 -29.810 ;
        RECT 1678.020 -29.820 1681.020 -29.810 ;
        RECT 1858.020 -29.820 1861.020 -29.810 ;
        RECT 2038.020 -29.820 2041.020 -29.810 ;
        RECT 2218.020 -29.820 2221.020 -29.810 ;
        RECT 2398.020 -29.820 2401.020 -29.810 ;
        RECT 2578.020 -29.820 2581.020 -29.810 ;
        RECT 2758.020 -29.820 2761.020 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 58.020 -32.830 61.020 -32.820 ;
        RECT 238.020 -32.830 241.020 -32.820 ;
        RECT 418.020 -32.830 421.020 -32.820 ;
        RECT 598.020 -32.830 601.020 -32.820 ;
        RECT 778.020 -32.830 781.020 -32.820 ;
        RECT 958.020 -32.830 961.020 -32.820 ;
        RECT 1138.020 -32.830 1141.020 -32.820 ;
        RECT 1318.020 -32.830 1321.020 -32.820 ;
        RECT 1498.020 -32.830 1501.020 -32.820 ;
        RECT 1678.020 -32.830 1681.020 -32.820 ;
        RECT 1858.020 -32.830 1861.020 -32.820 ;
        RECT 2038.020 -32.830 2041.020 -32.820 ;
        RECT 2218.020 -32.830 2221.020 -32.820 ;
        RECT 2398.020 -32.830 2401.020 -32.820 ;
        RECT 2578.020 -32.830 2581.020 -32.820 ;
        RECT 2758.020 -32.830 2761.020 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT 148.020 -37.520 151.020 3557.200 ;
        RECT 328.020 -37.520 331.020 3557.200 ;
        RECT 508.020 -37.520 511.020 3557.200 ;
        RECT 688.020 -37.520 691.020 3557.200 ;
        RECT 868.020 -37.520 871.020 3557.200 ;
        RECT 1048.020 -37.520 1051.020 3557.200 ;
        RECT 1228.020 -37.520 1231.020 3557.200 ;
        RECT 1408.020 -37.520 1411.020 3557.200 ;
        RECT 1588.020 -37.520 1591.020 3557.200 ;
        RECT 1768.020 -37.520 1771.020 3557.200 ;
        RECT 1948.020 -37.520 1951.020 3557.200 ;
        RECT 2128.020 -37.520 2131.020 3557.200 ;
        RECT 2308.020 -37.520 2311.020 3557.200 ;
        RECT 2488.020 -37.520 2491.020 3557.200 ;
        RECT 2668.020 -37.520 2671.020 3557.200 ;
        RECT 2848.020 -37.520 2851.020 3557.200 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT -41.970 3395.090 -40.790 3396.270 ;
        RECT -41.970 3393.490 -40.790 3394.670 ;
        RECT -41.970 3215.090 -40.790 3216.270 ;
        RECT -41.970 3213.490 -40.790 3214.670 ;
        RECT -41.970 3035.090 -40.790 3036.270 ;
        RECT -41.970 3033.490 -40.790 3034.670 ;
        RECT -41.970 2855.090 -40.790 2856.270 ;
        RECT -41.970 2853.490 -40.790 2854.670 ;
        RECT -41.970 2675.090 -40.790 2676.270 ;
        RECT -41.970 2673.490 -40.790 2674.670 ;
        RECT -41.970 2495.090 -40.790 2496.270 ;
        RECT -41.970 2493.490 -40.790 2494.670 ;
        RECT -41.970 2315.090 -40.790 2316.270 ;
        RECT -41.970 2313.490 -40.790 2314.670 ;
        RECT -41.970 2135.090 -40.790 2136.270 ;
        RECT -41.970 2133.490 -40.790 2134.670 ;
        RECT -41.970 1955.090 -40.790 1956.270 ;
        RECT -41.970 1953.490 -40.790 1954.670 ;
        RECT -41.970 1775.090 -40.790 1776.270 ;
        RECT -41.970 1773.490 -40.790 1774.670 ;
        RECT -41.970 1595.090 -40.790 1596.270 ;
        RECT -41.970 1593.490 -40.790 1594.670 ;
        RECT -41.970 1415.090 -40.790 1416.270 ;
        RECT -41.970 1413.490 -40.790 1414.670 ;
        RECT -41.970 1235.090 -40.790 1236.270 ;
        RECT -41.970 1233.490 -40.790 1234.670 ;
        RECT -41.970 1055.090 -40.790 1056.270 ;
        RECT -41.970 1053.490 -40.790 1054.670 ;
        RECT -41.970 875.090 -40.790 876.270 ;
        RECT -41.970 873.490 -40.790 874.670 ;
        RECT -41.970 695.090 -40.790 696.270 ;
        RECT -41.970 693.490 -40.790 694.670 ;
        RECT -41.970 515.090 -40.790 516.270 ;
        RECT -41.970 513.490 -40.790 514.670 ;
        RECT -41.970 335.090 -40.790 336.270 ;
        RECT -41.970 333.490 -40.790 334.670 ;
        RECT -41.970 155.090 -40.790 156.270 ;
        RECT -41.970 153.490 -40.790 154.670 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 148.930 3555.910 150.110 3557.090 ;
        RECT 148.930 3554.310 150.110 3555.490 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.810 150.110 -34.630 ;
        RECT 148.930 -37.410 150.110 -36.230 ;
        RECT 328.930 3555.910 330.110 3557.090 ;
        RECT 328.930 3554.310 330.110 3555.490 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 328.930 2675.090 330.110 2676.270 ;
        RECT 328.930 2673.490 330.110 2674.670 ;
        RECT 328.930 2495.090 330.110 2496.270 ;
        RECT 328.930 2493.490 330.110 2494.670 ;
        RECT 328.930 2315.090 330.110 2316.270 ;
        RECT 328.930 2313.490 330.110 2314.670 ;
        RECT 328.930 2135.090 330.110 2136.270 ;
        RECT 328.930 2133.490 330.110 2134.670 ;
        RECT 328.930 1955.090 330.110 1956.270 ;
        RECT 328.930 1953.490 330.110 1954.670 ;
        RECT 328.930 1775.090 330.110 1776.270 ;
        RECT 328.930 1773.490 330.110 1774.670 ;
        RECT 328.930 1595.090 330.110 1596.270 ;
        RECT 328.930 1593.490 330.110 1594.670 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.810 330.110 -34.630 ;
        RECT 328.930 -37.410 330.110 -36.230 ;
        RECT 508.930 3555.910 510.110 3557.090 ;
        RECT 508.930 3554.310 510.110 3555.490 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 508.930 3215.090 510.110 3216.270 ;
        RECT 508.930 3213.490 510.110 3214.670 ;
        RECT 508.930 3035.090 510.110 3036.270 ;
        RECT 508.930 3033.490 510.110 3034.670 ;
        RECT 508.930 2855.090 510.110 2856.270 ;
        RECT 508.930 2853.490 510.110 2854.670 ;
        RECT 508.930 2675.090 510.110 2676.270 ;
        RECT 508.930 2673.490 510.110 2674.670 ;
        RECT 508.930 2495.090 510.110 2496.270 ;
        RECT 508.930 2493.490 510.110 2494.670 ;
        RECT 508.930 2315.090 510.110 2316.270 ;
        RECT 508.930 2313.490 510.110 2314.670 ;
        RECT 508.930 2135.090 510.110 2136.270 ;
        RECT 508.930 2133.490 510.110 2134.670 ;
        RECT 508.930 1955.090 510.110 1956.270 ;
        RECT 508.930 1953.490 510.110 1954.670 ;
        RECT 508.930 1775.090 510.110 1776.270 ;
        RECT 508.930 1773.490 510.110 1774.670 ;
        RECT 508.930 1595.090 510.110 1596.270 ;
        RECT 508.930 1593.490 510.110 1594.670 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.810 510.110 -34.630 ;
        RECT 508.930 -37.410 510.110 -36.230 ;
        RECT 688.930 3555.910 690.110 3557.090 ;
        RECT 688.930 3554.310 690.110 3555.490 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 688.930 3215.090 690.110 3216.270 ;
        RECT 688.930 3213.490 690.110 3214.670 ;
        RECT 688.930 3035.090 690.110 3036.270 ;
        RECT 688.930 3033.490 690.110 3034.670 ;
        RECT 688.930 2855.090 690.110 2856.270 ;
        RECT 688.930 2853.490 690.110 2854.670 ;
        RECT 688.930 2675.090 690.110 2676.270 ;
        RECT 688.930 2673.490 690.110 2674.670 ;
        RECT 688.930 2495.090 690.110 2496.270 ;
        RECT 688.930 2493.490 690.110 2494.670 ;
        RECT 688.930 2315.090 690.110 2316.270 ;
        RECT 688.930 2313.490 690.110 2314.670 ;
        RECT 688.930 2135.090 690.110 2136.270 ;
        RECT 688.930 2133.490 690.110 2134.670 ;
        RECT 688.930 1955.090 690.110 1956.270 ;
        RECT 688.930 1953.490 690.110 1954.670 ;
        RECT 688.930 1775.090 690.110 1776.270 ;
        RECT 688.930 1773.490 690.110 1774.670 ;
        RECT 688.930 1595.090 690.110 1596.270 ;
        RECT 688.930 1593.490 690.110 1594.670 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 688.930 875.090 690.110 876.270 ;
        RECT 688.930 873.490 690.110 874.670 ;
        RECT 688.930 695.090 690.110 696.270 ;
        RECT 688.930 693.490 690.110 694.670 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.810 690.110 -34.630 ;
        RECT 688.930 -37.410 690.110 -36.230 ;
        RECT 868.930 3555.910 870.110 3557.090 ;
        RECT 868.930 3554.310 870.110 3555.490 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 868.930 2675.090 870.110 2676.270 ;
        RECT 868.930 2673.490 870.110 2674.670 ;
        RECT 868.930 2495.090 870.110 2496.270 ;
        RECT 868.930 2493.490 870.110 2494.670 ;
        RECT 868.930 2315.090 870.110 2316.270 ;
        RECT 868.930 2313.490 870.110 2314.670 ;
        RECT 868.930 2135.090 870.110 2136.270 ;
        RECT 868.930 2133.490 870.110 2134.670 ;
        RECT 868.930 1955.090 870.110 1956.270 ;
        RECT 868.930 1953.490 870.110 1954.670 ;
        RECT 868.930 1775.090 870.110 1776.270 ;
        RECT 868.930 1773.490 870.110 1774.670 ;
        RECT 868.930 1595.090 870.110 1596.270 ;
        RECT 868.930 1593.490 870.110 1594.670 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 868.930 875.090 870.110 876.270 ;
        RECT 868.930 873.490 870.110 874.670 ;
        RECT 868.930 695.090 870.110 696.270 ;
        RECT 868.930 693.490 870.110 694.670 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.810 870.110 -34.630 ;
        RECT 868.930 -37.410 870.110 -36.230 ;
        RECT 1048.930 3555.910 1050.110 3557.090 ;
        RECT 1048.930 3554.310 1050.110 3555.490 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1048.930 3215.090 1050.110 3216.270 ;
        RECT 1048.930 3213.490 1050.110 3214.670 ;
        RECT 1048.930 3035.090 1050.110 3036.270 ;
        RECT 1048.930 3033.490 1050.110 3034.670 ;
        RECT 1048.930 2855.090 1050.110 2856.270 ;
        RECT 1048.930 2853.490 1050.110 2854.670 ;
        RECT 1048.930 2675.090 1050.110 2676.270 ;
        RECT 1048.930 2673.490 1050.110 2674.670 ;
        RECT 1048.930 2495.090 1050.110 2496.270 ;
        RECT 1048.930 2493.490 1050.110 2494.670 ;
        RECT 1048.930 2315.090 1050.110 2316.270 ;
        RECT 1048.930 2313.490 1050.110 2314.670 ;
        RECT 1048.930 2135.090 1050.110 2136.270 ;
        RECT 1048.930 2133.490 1050.110 2134.670 ;
        RECT 1048.930 1955.090 1050.110 1956.270 ;
        RECT 1048.930 1953.490 1050.110 1954.670 ;
        RECT 1048.930 1775.090 1050.110 1776.270 ;
        RECT 1048.930 1773.490 1050.110 1774.670 ;
        RECT 1048.930 1595.090 1050.110 1596.270 ;
        RECT 1048.930 1593.490 1050.110 1594.670 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1048.930 875.090 1050.110 876.270 ;
        RECT 1048.930 873.490 1050.110 874.670 ;
        RECT 1048.930 695.090 1050.110 696.270 ;
        RECT 1048.930 693.490 1050.110 694.670 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.810 1050.110 -34.630 ;
        RECT 1048.930 -37.410 1050.110 -36.230 ;
        RECT 1228.930 3555.910 1230.110 3557.090 ;
        RECT 1228.930 3554.310 1230.110 3555.490 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1228.930 3215.090 1230.110 3216.270 ;
        RECT 1228.930 3213.490 1230.110 3214.670 ;
        RECT 1228.930 3035.090 1230.110 3036.270 ;
        RECT 1228.930 3033.490 1230.110 3034.670 ;
        RECT 1228.930 2855.090 1230.110 2856.270 ;
        RECT 1228.930 2853.490 1230.110 2854.670 ;
        RECT 1228.930 2675.090 1230.110 2676.270 ;
        RECT 1228.930 2673.490 1230.110 2674.670 ;
        RECT 1228.930 2495.090 1230.110 2496.270 ;
        RECT 1228.930 2493.490 1230.110 2494.670 ;
        RECT 1228.930 2315.090 1230.110 2316.270 ;
        RECT 1228.930 2313.490 1230.110 2314.670 ;
        RECT 1228.930 2135.090 1230.110 2136.270 ;
        RECT 1228.930 2133.490 1230.110 2134.670 ;
        RECT 1228.930 1955.090 1230.110 1956.270 ;
        RECT 1228.930 1953.490 1230.110 1954.670 ;
        RECT 1228.930 1775.090 1230.110 1776.270 ;
        RECT 1228.930 1773.490 1230.110 1774.670 ;
        RECT 1228.930 1595.090 1230.110 1596.270 ;
        RECT 1228.930 1593.490 1230.110 1594.670 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1228.930 875.090 1230.110 876.270 ;
        RECT 1228.930 873.490 1230.110 874.670 ;
        RECT 1228.930 695.090 1230.110 696.270 ;
        RECT 1228.930 693.490 1230.110 694.670 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.810 1230.110 -34.630 ;
        RECT 1228.930 -37.410 1230.110 -36.230 ;
        RECT 1408.930 3555.910 1410.110 3557.090 ;
        RECT 1408.930 3554.310 1410.110 3555.490 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1408.930 2675.090 1410.110 2676.270 ;
        RECT 1408.930 2673.490 1410.110 2674.670 ;
        RECT 1408.930 2495.090 1410.110 2496.270 ;
        RECT 1408.930 2493.490 1410.110 2494.670 ;
        RECT 1408.930 2315.090 1410.110 2316.270 ;
        RECT 1408.930 2313.490 1410.110 2314.670 ;
        RECT 1408.930 2135.090 1410.110 2136.270 ;
        RECT 1408.930 2133.490 1410.110 2134.670 ;
        RECT 1408.930 1955.090 1410.110 1956.270 ;
        RECT 1408.930 1953.490 1410.110 1954.670 ;
        RECT 1408.930 1775.090 1410.110 1776.270 ;
        RECT 1408.930 1773.490 1410.110 1774.670 ;
        RECT 1408.930 1595.090 1410.110 1596.270 ;
        RECT 1408.930 1593.490 1410.110 1594.670 ;
        RECT 1408.930 1415.090 1410.110 1416.270 ;
        RECT 1408.930 1413.490 1410.110 1414.670 ;
        RECT 1408.930 1235.090 1410.110 1236.270 ;
        RECT 1408.930 1233.490 1410.110 1234.670 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1408.930 875.090 1410.110 876.270 ;
        RECT 1408.930 873.490 1410.110 874.670 ;
        RECT 1408.930 695.090 1410.110 696.270 ;
        RECT 1408.930 693.490 1410.110 694.670 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.810 1410.110 -34.630 ;
        RECT 1408.930 -37.410 1410.110 -36.230 ;
        RECT 1588.930 3555.910 1590.110 3557.090 ;
        RECT 1588.930 3554.310 1590.110 3555.490 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1588.930 3035.090 1590.110 3036.270 ;
        RECT 1588.930 3033.490 1590.110 3034.670 ;
        RECT 1588.930 2855.090 1590.110 2856.270 ;
        RECT 1588.930 2853.490 1590.110 2854.670 ;
        RECT 1588.930 2675.090 1590.110 2676.270 ;
        RECT 1588.930 2673.490 1590.110 2674.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1588.930 2315.090 1590.110 2316.270 ;
        RECT 1588.930 2313.490 1590.110 2314.670 ;
        RECT 1588.930 2135.090 1590.110 2136.270 ;
        RECT 1588.930 2133.490 1590.110 2134.670 ;
        RECT 1588.930 1955.090 1590.110 1956.270 ;
        RECT 1588.930 1953.490 1590.110 1954.670 ;
        RECT 1588.930 1775.090 1590.110 1776.270 ;
        RECT 1588.930 1773.490 1590.110 1774.670 ;
        RECT 1588.930 1595.090 1590.110 1596.270 ;
        RECT 1588.930 1593.490 1590.110 1594.670 ;
        RECT 1588.930 1415.090 1590.110 1416.270 ;
        RECT 1588.930 1413.490 1590.110 1414.670 ;
        RECT 1588.930 1235.090 1590.110 1236.270 ;
        RECT 1588.930 1233.490 1590.110 1234.670 ;
        RECT 1588.930 1055.090 1590.110 1056.270 ;
        RECT 1588.930 1053.490 1590.110 1054.670 ;
        RECT 1588.930 875.090 1590.110 876.270 ;
        RECT 1588.930 873.490 1590.110 874.670 ;
        RECT 1588.930 695.090 1590.110 696.270 ;
        RECT 1588.930 693.490 1590.110 694.670 ;
        RECT 1588.930 515.090 1590.110 516.270 ;
        RECT 1588.930 513.490 1590.110 514.670 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.810 1590.110 -34.630 ;
        RECT 1588.930 -37.410 1590.110 -36.230 ;
        RECT 1768.930 3555.910 1770.110 3557.090 ;
        RECT 1768.930 3554.310 1770.110 3555.490 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1768.930 3035.090 1770.110 3036.270 ;
        RECT 1768.930 3033.490 1770.110 3034.670 ;
        RECT 1768.930 2855.090 1770.110 2856.270 ;
        RECT 1768.930 2853.490 1770.110 2854.670 ;
        RECT 1768.930 2675.090 1770.110 2676.270 ;
        RECT 1768.930 2673.490 1770.110 2674.670 ;
        RECT 1768.930 2495.090 1770.110 2496.270 ;
        RECT 1768.930 2493.490 1770.110 2494.670 ;
        RECT 1768.930 2315.090 1770.110 2316.270 ;
        RECT 1768.930 2313.490 1770.110 2314.670 ;
        RECT 1768.930 2135.090 1770.110 2136.270 ;
        RECT 1768.930 2133.490 1770.110 2134.670 ;
        RECT 1768.930 1955.090 1770.110 1956.270 ;
        RECT 1768.930 1953.490 1770.110 1954.670 ;
        RECT 1768.930 1775.090 1770.110 1776.270 ;
        RECT 1768.930 1773.490 1770.110 1774.670 ;
        RECT 1768.930 1595.090 1770.110 1596.270 ;
        RECT 1768.930 1593.490 1770.110 1594.670 ;
        RECT 1768.930 1415.090 1770.110 1416.270 ;
        RECT 1768.930 1413.490 1770.110 1414.670 ;
        RECT 1768.930 1235.090 1770.110 1236.270 ;
        RECT 1768.930 1233.490 1770.110 1234.670 ;
        RECT 1768.930 1055.090 1770.110 1056.270 ;
        RECT 1768.930 1053.490 1770.110 1054.670 ;
        RECT 1768.930 875.090 1770.110 876.270 ;
        RECT 1768.930 873.490 1770.110 874.670 ;
        RECT 1768.930 695.090 1770.110 696.270 ;
        RECT 1768.930 693.490 1770.110 694.670 ;
        RECT 1768.930 515.090 1770.110 516.270 ;
        RECT 1768.930 513.490 1770.110 514.670 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.810 1770.110 -34.630 ;
        RECT 1768.930 -37.410 1770.110 -36.230 ;
        RECT 1948.930 3555.910 1950.110 3557.090 ;
        RECT 1948.930 3554.310 1950.110 3555.490 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 1948.930 2855.090 1950.110 2856.270 ;
        RECT 1948.930 2853.490 1950.110 2854.670 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 1948.930 2495.090 1950.110 2496.270 ;
        RECT 1948.930 2493.490 1950.110 2494.670 ;
        RECT 1948.930 2315.090 1950.110 2316.270 ;
        RECT 1948.930 2313.490 1950.110 2314.670 ;
        RECT 1948.930 2135.090 1950.110 2136.270 ;
        RECT 1948.930 2133.490 1950.110 2134.670 ;
        RECT 1948.930 1955.090 1950.110 1956.270 ;
        RECT 1948.930 1953.490 1950.110 1954.670 ;
        RECT 1948.930 1775.090 1950.110 1776.270 ;
        RECT 1948.930 1773.490 1950.110 1774.670 ;
        RECT 1948.930 1595.090 1950.110 1596.270 ;
        RECT 1948.930 1593.490 1950.110 1594.670 ;
        RECT 1948.930 1415.090 1950.110 1416.270 ;
        RECT 1948.930 1413.490 1950.110 1414.670 ;
        RECT 1948.930 1235.090 1950.110 1236.270 ;
        RECT 1948.930 1233.490 1950.110 1234.670 ;
        RECT 1948.930 1055.090 1950.110 1056.270 ;
        RECT 1948.930 1053.490 1950.110 1054.670 ;
        RECT 1948.930 875.090 1950.110 876.270 ;
        RECT 1948.930 873.490 1950.110 874.670 ;
        RECT 1948.930 695.090 1950.110 696.270 ;
        RECT 1948.930 693.490 1950.110 694.670 ;
        RECT 1948.930 515.090 1950.110 516.270 ;
        RECT 1948.930 513.490 1950.110 514.670 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.810 1950.110 -34.630 ;
        RECT 1948.930 -37.410 1950.110 -36.230 ;
        RECT 2128.930 3555.910 2130.110 3557.090 ;
        RECT 2128.930 3554.310 2130.110 3555.490 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2128.930 2675.090 2130.110 2676.270 ;
        RECT 2128.930 2673.490 2130.110 2674.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2128.930 2315.090 2130.110 2316.270 ;
        RECT 2128.930 2313.490 2130.110 2314.670 ;
        RECT 2128.930 2135.090 2130.110 2136.270 ;
        RECT 2128.930 2133.490 2130.110 2134.670 ;
        RECT 2128.930 1955.090 2130.110 1956.270 ;
        RECT 2128.930 1953.490 2130.110 1954.670 ;
        RECT 2128.930 1775.090 2130.110 1776.270 ;
        RECT 2128.930 1773.490 2130.110 1774.670 ;
        RECT 2128.930 1595.090 2130.110 1596.270 ;
        RECT 2128.930 1593.490 2130.110 1594.670 ;
        RECT 2128.930 1415.090 2130.110 1416.270 ;
        RECT 2128.930 1413.490 2130.110 1414.670 ;
        RECT 2128.930 1235.090 2130.110 1236.270 ;
        RECT 2128.930 1233.490 2130.110 1234.670 ;
        RECT 2128.930 1055.090 2130.110 1056.270 ;
        RECT 2128.930 1053.490 2130.110 1054.670 ;
        RECT 2128.930 875.090 2130.110 876.270 ;
        RECT 2128.930 873.490 2130.110 874.670 ;
        RECT 2128.930 695.090 2130.110 696.270 ;
        RECT 2128.930 693.490 2130.110 694.670 ;
        RECT 2128.930 515.090 2130.110 516.270 ;
        RECT 2128.930 513.490 2130.110 514.670 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.810 2130.110 -34.630 ;
        RECT 2128.930 -37.410 2130.110 -36.230 ;
        RECT 2308.930 3555.910 2310.110 3557.090 ;
        RECT 2308.930 3554.310 2310.110 3555.490 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2308.930 3035.090 2310.110 3036.270 ;
        RECT 2308.930 3033.490 2310.110 3034.670 ;
        RECT 2308.930 2855.090 2310.110 2856.270 ;
        RECT 2308.930 2853.490 2310.110 2854.670 ;
        RECT 2308.930 2675.090 2310.110 2676.270 ;
        RECT 2308.930 2673.490 2310.110 2674.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2308.930 2315.090 2310.110 2316.270 ;
        RECT 2308.930 2313.490 2310.110 2314.670 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2308.930 1955.090 2310.110 1956.270 ;
        RECT 2308.930 1953.490 2310.110 1954.670 ;
        RECT 2308.930 1775.090 2310.110 1776.270 ;
        RECT 2308.930 1773.490 2310.110 1774.670 ;
        RECT 2308.930 1595.090 2310.110 1596.270 ;
        RECT 2308.930 1593.490 2310.110 1594.670 ;
        RECT 2308.930 1415.090 2310.110 1416.270 ;
        RECT 2308.930 1413.490 2310.110 1414.670 ;
        RECT 2308.930 1235.090 2310.110 1236.270 ;
        RECT 2308.930 1233.490 2310.110 1234.670 ;
        RECT 2308.930 1055.090 2310.110 1056.270 ;
        RECT 2308.930 1053.490 2310.110 1054.670 ;
        RECT 2308.930 875.090 2310.110 876.270 ;
        RECT 2308.930 873.490 2310.110 874.670 ;
        RECT 2308.930 695.090 2310.110 696.270 ;
        RECT 2308.930 693.490 2310.110 694.670 ;
        RECT 2308.930 515.090 2310.110 516.270 ;
        RECT 2308.930 513.490 2310.110 514.670 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.810 2310.110 -34.630 ;
        RECT 2308.930 -37.410 2310.110 -36.230 ;
        RECT 2488.930 3555.910 2490.110 3557.090 ;
        RECT 2488.930 3554.310 2490.110 3555.490 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2488.930 3035.090 2490.110 3036.270 ;
        RECT 2488.930 3033.490 2490.110 3034.670 ;
        RECT 2488.930 2855.090 2490.110 2856.270 ;
        RECT 2488.930 2853.490 2490.110 2854.670 ;
        RECT 2488.930 2675.090 2490.110 2676.270 ;
        RECT 2488.930 2673.490 2490.110 2674.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2488.930 2315.090 2490.110 2316.270 ;
        RECT 2488.930 2313.490 2490.110 2314.670 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2488.930 1955.090 2490.110 1956.270 ;
        RECT 2488.930 1953.490 2490.110 1954.670 ;
        RECT 2488.930 1775.090 2490.110 1776.270 ;
        RECT 2488.930 1773.490 2490.110 1774.670 ;
        RECT 2488.930 1595.090 2490.110 1596.270 ;
        RECT 2488.930 1593.490 2490.110 1594.670 ;
        RECT 2488.930 1415.090 2490.110 1416.270 ;
        RECT 2488.930 1413.490 2490.110 1414.670 ;
        RECT 2488.930 1235.090 2490.110 1236.270 ;
        RECT 2488.930 1233.490 2490.110 1234.670 ;
        RECT 2488.930 1055.090 2490.110 1056.270 ;
        RECT 2488.930 1053.490 2490.110 1054.670 ;
        RECT 2488.930 875.090 2490.110 876.270 ;
        RECT 2488.930 873.490 2490.110 874.670 ;
        RECT 2488.930 695.090 2490.110 696.270 ;
        RECT 2488.930 693.490 2490.110 694.670 ;
        RECT 2488.930 515.090 2490.110 516.270 ;
        RECT 2488.930 513.490 2490.110 514.670 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.810 2490.110 -34.630 ;
        RECT 2488.930 -37.410 2490.110 -36.230 ;
        RECT 2668.930 3555.910 2670.110 3557.090 ;
        RECT 2668.930 3554.310 2670.110 3555.490 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.810 2670.110 -34.630 ;
        RECT 2668.930 -37.410 2670.110 -36.230 ;
        RECT 2848.930 3555.910 2850.110 3557.090 ;
        RECT 2848.930 3554.310 2850.110 3555.490 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.810 2850.110 -34.630 ;
        RECT 2848.930 -37.410 2850.110 -36.230 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT 2960.410 3395.090 2961.590 3396.270 ;
        RECT 2960.410 3393.490 2961.590 3394.670 ;
        RECT 2960.410 3215.090 2961.590 3216.270 ;
        RECT 2960.410 3213.490 2961.590 3214.670 ;
        RECT 2960.410 3035.090 2961.590 3036.270 ;
        RECT 2960.410 3033.490 2961.590 3034.670 ;
        RECT 2960.410 2855.090 2961.590 2856.270 ;
        RECT 2960.410 2853.490 2961.590 2854.670 ;
        RECT 2960.410 2675.090 2961.590 2676.270 ;
        RECT 2960.410 2673.490 2961.590 2674.670 ;
        RECT 2960.410 2495.090 2961.590 2496.270 ;
        RECT 2960.410 2493.490 2961.590 2494.670 ;
        RECT 2960.410 2315.090 2961.590 2316.270 ;
        RECT 2960.410 2313.490 2961.590 2314.670 ;
        RECT 2960.410 2135.090 2961.590 2136.270 ;
        RECT 2960.410 2133.490 2961.590 2134.670 ;
        RECT 2960.410 1955.090 2961.590 1956.270 ;
        RECT 2960.410 1953.490 2961.590 1954.670 ;
        RECT 2960.410 1775.090 2961.590 1776.270 ;
        RECT 2960.410 1773.490 2961.590 1774.670 ;
        RECT 2960.410 1595.090 2961.590 1596.270 ;
        RECT 2960.410 1593.490 2961.590 1594.670 ;
        RECT 2960.410 1415.090 2961.590 1416.270 ;
        RECT 2960.410 1413.490 2961.590 1414.670 ;
        RECT 2960.410 1235.090 2961.590 1236.270 ;
        RECT 2960.410 1233.490 2961.590 1234.670 ;
        RECT 2960.410 1055.090 2961.590 1056.270 ;
        RECT 2960.410 1053.490 2961.590 1054.670 ;
        RECT 2960.410 875.090 2961.590 876.270 ;
        RECT 2960.410 873.490 2961.590 874.670 ;
        RECT 2960.410 695.090 2961.590 696.270 ;
        RECT 2960.410 693.490 2961.590 694.670 ;
        RECT 2960.410 515.090 2961.590 516.270 ;
        RECT 2960.410 513.490 2961.590 514.670 ;
        RECT 2960.410 335.090 2961.590 336.270 ;
        RECT 2960.410 333.490 2961.590 334.670 ;
        RECT 2960.410 155.090 2961.590 156.270 ;
        RECT 2960.410 153.490 2961.590 154.670 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 148.020 3557.200 151.020 3557.210 ;
        RECT 328.020 3557.200 331.020 3557.210 ;
        RECT 508.020 3557.200 511.020 3557.210 ;
        RECT 688.020 3557.200 691.020 3557.210 ;
        RECT 868.020 3557.200 871.020 3557.210 ;
        RECT 1048.020 3557.200 1051.020 3557.210 ;
        RECT 1228.020 3557.200 1231.020 3557.210 ;
        RECT 1408.020 3557.200 1411.020 3557.210 ;
        RECT 1588.020 3557.200 1591.020 3557.210 ;
        RECT 1768.020 3557.200 1771.020 3557.210 ;
        RECT 1948.020 3557.200 1951.020 3557.210 ;
        RECT 2128.020 3557.200 2131.020 3557.210 ;
        RECT 2308.020 3557.200 2311.020 3557.210 ;
        RECT 2488.020 3557.200 2491.020 3557.210 ;
        RECT 2668.020 3557.200 2671.020 3557.210 ;
        RECT 2848.020 3557.200 2851.020 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 148.020 3554.190 151.020 3554.200 ;
        RECT 328.020 3554.190 331.020 3554.200 ;
        RECT 508.020 3554.190 511.020 3554.200 ;
        RECT 688.020 3554.190 691.020 3554.200 ;
        RECT 868.020 3554.190 871.020 3554.200 ;
        RECT 1048.020 3554.190 1051.020 3554.200 ;
        RECT 1228.020 3554.190 1231.020 3554.200 ;
        RECT 1408.020 3554.190 1411.020 3554.200 ;
        RECT 1588.020 3554.190 1591.020 3554.200 ;
        RECT 1768.020 3554.190 1771.020 3554.200 ;
        RECT 1948.020 3554.190 1951.020 3554.200 ;
        RECT 2128.020 3554.190 2131.020 3554.200 ;
        RECT 2308.020 3554.190 2311.020 3554.200 ;
        RECT 2488.020 3554.190 2491.020 3554.200 ;
        RECT 2668.020 3554.190 2671.020 3554.200 ;
        RECT 2848.020 3554.190 2851.020 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -42.880 3396.380 -39.880 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2959.500 3396.380 2962.500 3396.390 ;
        RECT -42.880 3393.380 2962.500 3396.380 ;
        RECT -42.880 3393.370 -39.880 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2959.500 3393.370 2962.500 3393.380 ;
        RECT -42.880 3216.380 -39.880 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 508.020 3216.380 511.020 3216.390 ;
        RECT 688.020 3216.380 691.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1048.020 3216.380 1051.020 3216.390 ;
        RECT 1228.020 3216.380 1231.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2959.500 3216.380 2962.500 3216.390 ;
        RECT -42.880 3213.380 2962.500 3216.380 ;
        RECT -42.880 3213.370 -39.880 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 508.020 3213.370 511.020 3213.380 ;
        RECT 688.020 3213.370 691.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1048.020 3213.370 1051.020 3213.380 ;
        RECT 1228.020 3213.370 1231.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2959.500 3213.370 2962.500 3213.380 ;
        RECT -42.880 3036.380 -39.880 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 508.020 3036.380 511.020 3036.390 ;
        RECT 688.020 3036.380 691.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1048.020 3036.380 1051.020 3036.390 ;
        RECT 1228.020 3036.380 1231.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1588.020 3036.380 1591.020 3036.390 ;
        RECT 1768.020 3036.380 1771.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2308.020 3036.380 2311.020 3036.390 ;
        RECT 2488.020 3036.380 2491.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2959.500 3036.380 2962.500 3036.390 ;
        RECT -42.880 3033.380 2962.500 3036.380 ;
        RECT -42.880 3033.370 -39.880 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 508.020 3033.370 511.020 3033.380 ;
        RECT 688.020 3033.370 691.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1048.020 3033.370 1051.020 3033.380 ;
        RECT 1228.020 3033.370 1231.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1588.020 3033.370 1591.020 3033.380 ;
        RECT 1768.020 3033.370 1771.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2308.020 3033.370 2311.020 3033.380 ;
        RECT 2488.020 3033.370 2491.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2959.500 3033.370 2962.500 3033.380 ;
        RECT -42.880 2856.380 -39.880 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 508.020 2856.380 511.020 2856.390 ;
        RECT 688.020 2856.380 691.020 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1048.020 2856.380 1051.020 2856.390 ;
        RECT 1228.020 2856.380 1231.020 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1588.020 2856.380 1591.020 2856.390 ;
        RECT 1768.020 2856.380 1771.020 2856.390 ;
        RECT 1948.020 2856.380 1951.020 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2308.020 2856.380 2311.020 2856.390 ;
        RECT 2488.020 2856.380 2491.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2959.500 2856.380 2962.500 2856.390 ;
        RECT -42.880 2853.380 2962.500 2856.380 ;
        RECT -42.880 2853.370 -39.880 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 508.020 2853.370 511.020 2853.380 ;
        RECT 688.020 2853.370 691.020 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1048.020 2853.370 1051.020 2853.380 ;
        RECT 1228.020 2853.370 1231.020 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1588.020 2853.370 1591.020 2853.380 ;
        RECT 1768.020 2853.370 1771.020 2853.380 ;
        RECT 1948.020 2853.370 1951.020 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2308.020 2853.370 2311.020 2853.380 ;
        RECT 2488.020 2853.370 2491.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2959.500 2853.370 2962.500 2853.380 ;
        RECT -42.880 2676.380 -39.880 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 328.020 2676.380 331.020 2676.390 ;
        RECT 508.020 2676.380 511.020 2676.390 ;
        RECT 688.020 2676.380 691.020 2676.390 ;
        RECT 868.020 2676.380 871.020 2676.390 ;
        RECT 1048.020 2676.380 1051.020 2676.390 ;
        RECT 1228.020 2676.380 1231.020 2676.390 ;
        RECT 1408.020 2676.380 1411.020 2676.390 ;
        RECT 1588.020 2676.380 1591.020 2676.390 ;
        RECT 1768.020 2676.380 1771.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2128.020 2676.380 2131.020 2676.390 ;
        RECT 2308.020 2676.380 2311.020 2676.390 ;
        RECT 2488.020 2676.380 2491.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2959.500 2676.380 2962.500 2676.390 ;
        RECT -42.880 2673.380 2962.500 2676.380 ;
        RECT -42.880 2673.370 -39.880 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 328.020 2673.370 331.020 2673.380 ;
        RECT 508.020 2673.370 511.020 2673.380 ;
        RECT 688.020 2673.370 691.020 2673.380 ;
        RECT 868.020 2673.370 871.020 2673.380 ;
        RECT 1048.020 2673.370 1051.020 2673.380 ;
        RECT 1228.020 2673.370 1231.020 2673.380 ;
        RECT 1408.020 2673.370 1411.020 2673.380 ;
        RECT 1588.020 2673.370 1591.020 2673.380 ;
        RECT 1768.020 2673.370 1771.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2128.020 2673.370 2131.020 2673.380 ;
        RECT 2308.020 2673.370 2311.020 2673.380 ;
        RECT 2488.020 2673.370 2491.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2959.500 2673.370 2962.500 2673.380 ;
        RECT -42.880 2496.380 -39.880 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 328.020 2496.380 331.020 2496.390 ;
        RECT 508.020 2496.380 511.020 2496.390 ;
        RECT 688.020 2496.380 691.020 2496.390 ;
        RECT 868.020 2496.380 871.020 2496.390 ;
        RECT 1048.020 2496.380 1051.020 2496.390 ;
        RECT 1228.020 2496.380 1231.020 2496.390 ;
        RECT 1408.020 2496.380 1411.020 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 1768.020 2496.380 1771.020 2496.390 ;
        RECT 1948.020 2496.380 1951.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2959.500 2496.380 2962.500 2496.390 ;
        RECT -42.880 2493.380 2962.500 2496.380 ;
        RECT -42.880 2493.370 -39.880 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 328.020 2493.370 331.020 2493.380 ;
        RECT 508.020 2493.370 511.020 2493.380 ;
        RECT 688.020 2493.370 691.020 2493.380 ;
        RECT 868.020 2493.370 871.020 2493.380 ;
        RECT 1048.020 2493.370 1051.020 2493.380 ;
        RECT 1228.020 2493.370 1231.020 2493.380 ;
        RECT 1408.020 2493.370 1411.020 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 1768.020 2493.370 1771.020 2493.380 ;
        RECT 1948.020 2493.370 1951.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2959.500 2493.370 2962.500 2493.380 ;
        RECT -42.880 2316.380 -39.880 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 328.020 2316.380 331.020 2316.390 ;
        RECT 508.020 2316.380 511.020 2316.390 ;
        RECT 688.020 2316.380 691.020 2316.390 ;
        RECT 868.020 2316.380 871.020 2316.390 ;
        RECT 1048.020 2316.380 1051.020 2316.390 ;
        RECT 1228.020 2316.380 1231.020 2316.390 ;
        RECT 1408.020 2316.380 1411.020 2316.390 ;
        RECT 1588.020 2316.380 1591.020 2316.390 ;
        RECT 1768.020 2316.380 1771.020 2316.390 ;
        RECT 1948.020 2316.380 1951.020 2316.390 ;
        RECT 2128.020 2316.380 2131.020 2316.390 ;
        RECT 2308.020 2316.380 2311.020 2316.390 ;
        RECT 2488.020 2316.380 2491.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2959.500 2316.380 2962.500 2316.390 ;
        RECT -42.880 2313.380 2962.500 2316.380 ;
        RECT -42.880 2313.370 -39.880 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 328.020 2313.370 331.020 2313.380 ;
        RECT 508.020 2313.370 511.020 2313.380 ;
        RECT 688.020 2313.370 691.020 2313.380 ;
        RECT 868.020 2313.370 871.020 2313.380 ;
        RECT 1048.020 2313.370 1051.020 2313.380 ;
        RECT 1228.020 2313.370 1231.020 2313.380 ;
        RECT 1408.020 2313.370 1411.020 2313.380 ;
        RECT 1588.020 2313.370 1591.020 2313.380 ;
        RECT 1768.020 2313.370 1771.020 2313.380 ;
        RECT 1948.020 2313.370 1951.020 2313.380 ;
        RECT 2128.020 2313.370 2131.020 2313.380 ;
        RECT 2308.020 2313.370 2311.020 2313.380 ;
        RECT 2488.020 2313.370 2491.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2959.500 2313.370 2962.500 2313.380 ;
        RECT -42.880 2136.380 -39.880 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 328.020 2136.380 331.020 2136.390 ;
        RECT 508.020 2136.380 511.020 2136.390 ;
        RECT 688.020 2136.380 691.020 2136.390 ;
        RECT 868.020 2136.380 871.020 2136.390 ;
        RECT 1048.020 2136.380 1051.020 2136.390 ;
        RECT 1228.020 2136.380 1231.020 2136.390 ;
        RECT 1408.020 2136.380 1411.020 2136.390 ;
        RECT 1588.020 2136.380 1591.020 2136.390 ;
        RECT 1768.020 2136.380 1771.020 2136.390 ;
        RECT 1948.020 2136.380 1951.020 2136.390 ;
        RECT 2128.020 2136.380 2131.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2959.500 2136.380 2962.500 2136.390 ;
        RECT -42.880 2133.380 2962.500 2136.380 ;
        RECT -42.880 2133.370 -39.880 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 328.020 2133.370 331.020 2133.380 ;
        RECT 508.020 2133.370 511.020 2133.380 ;
        RECT 688.020 2133.370 691.020 2133.380 ;
        RECT 868.020 2133.370 871.020 2133.380 ;
        RECT 1048.020 2133.370 1051.020 2133.380 ;
        RECT 1228.020 2133.370 1231.020 2133.380 ;
        RECT 1408.020 2133.370 1411.020 2133.380 ;
        RECT 1588.020 2133.370 1591.020 2133.380 ;
        RECT 1768.020 2133.370 1771.020 2133.380 ;
        RECT 1948.020 2133.370 1951.020 2133.380 ;
        RECT 2128.020 2133.370 2131.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2959.500 2133.370 2962.500 2133.380 ;
        RECT -42.880 1956.380 -39.880 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 328.020 1956.380 331.020 1956.390 ;
        RECT 508.020 1956.380 511.020 1956.390 ;
        RECT 688.020 1956.380 691.020 1956.390 ;
        RECT 868.020 1956.380 871.020 1956.390 ;
        RECT 1048.020 1956.380 1051.020 1956.390 ;
        RECT 1228.020 1956.380 1231.020 1956.390 ;
        RECT 1408.020 1956.380 1411.020 1956.390 ;
        RECT 1588.020 1956.380 1591.020 1956.390 ;
        RECT 1768.020 1956.380 1771.020 1956.390 ;
        RECT 1948.020 1956.380 1951.020 1956.390 ;
        RECT 2128.020 1956.380 2131.020 1956.390 ;
        RECT 2308.020 1956.380 2311.020 1956.390 ;
        RECT 2488.020 1956.380 2491.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2959.500 1956.380 2962.500 1956.390 ;
        RECT -42.880 1953.380 2962.500 1956.380 ;
        RECT -42.880 1953.370 -39.880 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 328.020 1953.370 331.020 1953.380 ;
        RECT 508.020 1953.370 511.020 1953.380 ;
        RECT 688.020 1953.370 691.020 1953.380 ;
        RECT 868.020 1953.370 871.020 1953.380 ;
        RECT 1048.020 1953.370 1051.020 1953.380 ;
        RECT 1228.020 1953.370 1231.020 1953.380 ;
        RECT 1408.020 1953.370 1411.020 1953.380 ;
        RECT 1588.020 1953.370 1591.020 1953.380 ;
        RECT 1768.020 1953.370 1771.020 1953.380 ;
        RECT 1948.020 1953.370 1951.020 1953.380 ;
        RECT 2128.020 1953.370 2131.020 1953.380 ;
        RECT 2308.020 1953.370 2311.020 1953.380 ;
        RECT 2488.020 1953.370 2491.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2959.500 1953.370 2962.500 1953.380 ;
        RECT -42.880 1776.380 -39.880 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 328.020 1776.380 331.020 1776.390 ;
        RECT 508.020 1776.380 511.020 1776.390 ;
        RECT 688.020 1776.380 691.020 1776.390 ;
        RECT 868.020 1776.380 871.020 1776.390 ;
        RECT 1048.020 1776.380 1051.020 1776.390 ;
        RECT 1228.020 1776.380 1231.020 1776.390 ;
        RECT 1408.020 1776.380 1411.020 1776.390 ;
        RECT 1588.020 1776.380 1591.020 1776.390 ;
        RECT 1768.020 1776.380 1771.020 1776.390 ;
        RECT 1948.020 1776.380 1951.020 1776.390 ;
        RECT 2128.020 1776.380 2131.020 1776.390 ;
        RECT 2308.020 1776.380 2311.020 1776.390 ;
        RECT 2488.020 1776.380 2491.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2959.500 1776.380 2962.500 1776.390 ;
        RECT -42.880 1773.380 2962.500 1776.380 ;
        RECT -42.880 1773.370 -39.880 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 328.020 1773.370 331.020 1773.380 ;
        RECT 508.020 1773.370 511.020 1773.380 ;
        RECT 688.020 1773.370 691.020 1773.380 ;
        RECT 868.020 1773.370 871.020 1773.380 ;
        RECT 1048.020 1773.370 1051.020 1773.380 ;
        RECT 1228.020 1773.370 1231.020 1773.380 ;
        RECT 1408.020 1773.370 1411.020 1773.380 ;
        RECT 1588.020 1773.370 1591.020 1773.380 ;
        RECT 1768.020 1773.370 1771.020 1773.380 ;
        RECT 1948.020 1773.370 1951.020 1773.380 ;
        RECT 2128.020 1773.370 2131.020 1773.380 ;
        RECT 2308.020 1773.370 2311.020 1773.380 ;
        RECT 2488.020 1773.370 2491.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2959.500 1773.370 2962.500 1773.380 ;
        RECT -42.880 1596.380 -39.880 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 328.020 1596.380 331.020 1596.390 ;
        RECT 508.020 1596.380 511.020 1596.390 ;
        RECT 688.020 1596.380 691.020 1596.390 ;
        RECT 868.020 1596.380 871.020 1596.390 ;
        RECT 1048.020 1596.380 1051.020 1596.390 ;
        RECT 1228.020 1596.380 1231.020 1596.390 ;
        RECT 1408.020 1596.380 1411.020 1596.390 ;
        RECT 1588.020 1596.380 1591.020 1596.390 ;
        RECT 1768.020 1596.380 1771.020 1596.390 ;
        RECT 1948.020 1596.380 1951.020 1596.390 ;
        RECT 2128.020 1596.380 2131.020 1596.390 ;
        RECT 2308.020 1596.380 2311.020 1596.390 ;
        RECT 2488.020 1596.380 2491.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2959.500 1596.380 2962.500 1596.390 ;
        RECT -42.880 1593.380 2962.500 1596.380 ;
        RECT -42.880 1593.370 -39.880 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 328.020 1593.370 331.020 1593.380 ;
        RECT 508.020 1593.370 511.020 1593.380 ;
        RECT 688.020 1593.370 691.020 1593.380 ;
        RECT 868.020 1593.370 871.020 1593.380 ;
        RECT 1048.020 1593.370 1051.020 1593.380 ;
        RECT 1228.020 1593.370 1231.020 1593.380 ;
        RECT 1408.020 1593.370 1411.020 1593.380 ;
        RECT 1588.020 1593.370 1591.020 1593.380 ;
        RECT 1768.020 1593.370 1771.020 1593.380 ;
        RECT 1948.020 1593.370 1951.020 1593.380 ;
        RECT 2128.020 1593.370 2131.020 1593.380 ;
        RECT 2308.020 1593.370 2311.020 1593.380 ;
        RECT 2488.020 1593.370 2491.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2959.500 1593.370 2962.500 1593.380 ;
        RECT -42.880 1416.380 -39.880 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 1408.020 1416.380 1411.020 1416.390 ;
        RECT 1588.020 1416.380 1591.020 1416.390 ;
        RECT 1768.020 1416.380 1771.020 1416.390 ;
        RECT 1948.020 1416.380 1951.020 1416.390 ;
        RECT 2128.020 1416.380 2131.020 1416.390 ;
        RECT 2308.020 1416.380 2311.020 1416.390 ;
        RECT 2488.020 1416.380 2491.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2959.500 1416.380 2962.500 1416.390 ;
        RECT -42.880 1413.380 2962.500 1416.380 ;
        RECT -42.880 1413.370 -39.880 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 1408.020 1413.370 1411.020 1413.380 ;
        RECT 1588.020 1413.370 1591.020 1413.380 ;
        RECT 1768.020 1413.370 1771.020 1413.380 ;
        RECT 1948.020 1413.370 1951.020 1413.380 ;
        RECT 2128.020 1413.370 2131.020 1413.380 ;
        RECT 2308.020 1413.370 2311.020 1413.380 ;
        RECT 2488.020 1413.370 2491.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2959.500 1413.370 2962.500 1413.380 ;
        RECT -42.880 1236.380 -39.880 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 1408.020 1236.380 1411.020 1236.390 ;
        RECT 1588.020 1236.380 1591.020 1236.390 ;
        RECT 1768.020 1236.380 1771.020 1236.390 ;
        RECT 1948.020 1236.380 1951.020 1236.390 ;
        RECT 2128.020 1236.380 2131.020 1236.390 ;
        RECT 2308.020 1236.380 2311.020 1236.390 ;
        RECT 2488.020 1236.380 2491.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2959.500 1236.380 2962.500 1236.390 ;
        RECT -42.880 1233.380 2962.500 1236.380 ;
        RECT -42.880 1233.370 -39.880 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 1408.020 1233.370 1411.020 1233.380 ;
        RECT 1588.020 1233.370 1591.020 1233.380 ;
        RECT 1768.020 1233.370 1771.020 1233.380 ;
        RECT 1948.020 1233.370 1951.020 1233.380 ;
        RECT 2128.020 1233.370 2131.020 1233.380 ;
        RECT 2308.020 1233.370 2311.020 1233.380 ;
        RECT 2488.020 1233.370 2491.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2959.500 1233.370 2962.500 1233.380 ;
        RECT -42.880 1056.380 -39.880 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1588.020 1056.380 1591.020 1056.390 ;
        RECT 1768.020 1056.380 1771.020 1056.390 ;
        RECT 1948.020 1056.380 1951.020 1056.390 ;
        RECT 2128.020 1056.380 2131.020 1056.390 ;
        RECT 2308.020 1056.380 2311.020 1056.390 ;
        RECT 2488.020 1056.380 2491.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2959.500 1056.380 2962.500 1056.390 ;
        RECT -42.880 1053.380 2962.500 1056.380 ;
        RECT -42.880 1053.370 -39.880 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1588.020 1053.370 1591.020 1053.380 ;
        RECT 1768.020 1053.370 1771.020 1053.380 ;
        RECT 1948.020 1053.370 1951.020 1053.380 ;
        RECT 2128.020 1053.370 2131.020 1053.380 ;
        RECT 2308.020 1053.370 2311.020 1053.380 ;
        RECT 2488.020 1053.370 2491.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2959.500 1053.370 2962.500 1053.380 ;
        RECT -42.880 876.380 -39.880 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 688.020 876.380 691.020 876.390 ;
        RECT 868.020 876.380 871.020 876.390 ;
        RECT 1048.020 876.380 1051.020 876.390 ;
        RECT 1228.020 876.380 1231.020 876.390 ;
        RECT 1408.020 876.380 1411.020 876.390 ;
        RECT 1588.020 876.380 1591.020 876.390 ;
        RECT 1768.020 876.380 1771.020 876.390 ;
        RECT 1948.020 876.380 1951.020 876.390 ;
        RECT 2128.020 876.380 2131.020 876.390 ;
        RECT 2308.020 876.380 2311.020 876.390 ;
        RECT 2488.020 876.380 2491.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2959.500 876.380 2962.500 876.390 ;
        RECT -42.880 873.380 2962.500 876.380 ;
        RECT -42.880 873.370 -39.880 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 688.020 873.370 691.020 873.380 ;
        RECT 868.020 873.370 871.020 873.380 ;
        RECT 1048.020 873.370 1051.020 873.380 ;
        RECT 1228.020 873.370 1231.020 873.380 ;
        RECT 1408.020 873.370 1411.020 873.380 ;
        RECT 1588.020 873.370 1591.020 873.380 ;
        RECT 1768.020 873.370 1771.020 873.380 ;
        RECT 1948.020 873.370 1951.020 873.380 ;
        RECT 2128.020 873.370 2131.020 873.380 ;
        RECT 2308.020 873.370 2311.020 873.380 ;
        RECT 2488.020 873.370 2491.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2959.500 873.370 2962.500 873.380 ;
        RECT -42.880 696.380 -39.880 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 688.020 696.380 691.020 696.390 ;
        RECT 868.020 696.380 871.020 696.390 ;
        RECT 1048.020 696.380 1051.020 696.390 ;
        RECT 1228.020 696.380 1231.020 696.390 ;
        RECT 1408.020 696.380 1411.020 696.390 ;
        RECT 1588.020 696.380 1591.020 696.390 ;
        RECT 1768.020 696.380 1771.020 696.390 ;
        RECT 1948.020 696.380 1951.020 696.390 ;
        RECT 2128.020 696.380 2131.020 696.390 ;
        RECT 2308.020 696.380 2311.020 696.390 ;
        RECT 2488.020 696.380 2491.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2959.500 696.380 2962.500 696.390 ;
        RECT -42.880 693.380 2962.500 696.380 ;
        RECT -42.880 693.370 -39.880 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 688.020 693.370 691.020 693.380 ;
        RECT 868.020 693.370 871.020 693.380 ;
        RECT 1048.020 693.370 1051.020 693.380 ;
        RECT 1228.020 693.370 1231.020 693.380 ;
        RECT 1408.020 693.370 1411.020 693.380 ;
        RECT 1588.020 693.370 1591.020 693.380 ;
        RECT 1768.020 693.370 1771.020 693.380 ;
        RECT 1948.020 693.370 1951.020 693.380 ;
        RECT 2128.020 693.370 2131.020 693.380 ;
        RECT 2308.020 693.370 2311.020 693.380 ;
        RECT 2488.020 693.370 2491.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2959.500 693.370 2962.500 693.380 ;
        RECT -42.880 516.380 -39.880 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1588.020 516.380 1591.020 516.390 ;
        RECT 1768.020 516.380 1771.020 516.390 ;
        RECT 1948.020 516.380 1951.020 516.390 ;
        RECT 2128.020 516.380 2131.020 516.390 ;
        RECT 2308.020 516.380 2311.020 516.390 ;
        RECT 2488.020 516.380 2491.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2959.500 516.380 2962.500 516.390 ;
        RECT -42.880 513.380 2962.500 516.380 ;
        RECT -42.880 513.370 -39.880 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1588.020 513.370 1591.020 513.380 ;
        RECT 1768.020 513.370 1771.020 513.380 ;
        RECT 1948.020 513.370 1951.020 513.380 ;
        RECT 2128.020 513.370 2131.020 513.380 ;
        RECT 2308.020 513.370 2311.020 513.380 ;
        RECT 2488.020 513.370 2491.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2959.500 513.370 2962.500 513.380 ;
        RECT -42.880 336.380 -39.880 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2959.500 336.380 2962.500 336.390 ;
        RECT -42.880 333.380 2962.500 336.380 ;
        RECT -42.880 333.370 -39.880 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2959.500 333.370 2962.500 333.380 ;
        RECT -42.880 156.380 -39.880 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2959.500 156.380 2962.500 156.390 ;
        RECT -42.880 153.380 2962.500 156.380 ;
        RECT -42.880 153.370 -39.880 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2959.500 153.370 2962.500 153.380 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 148.020 -34.520 151.020 -34.510 ;
        RECT 328.020 -34.520 331.020 -34.510 ;
        RECT 508.020 -34.520 511.020 -34.510 ;
        RECT 688.020 -34.520 691.020 -34.510 ;
        RECT 868.020 -34.520 871.020 -34.510 ;
        RECT 1048.020 -34.520 1051.020 -34.510 ;
        RECT 1228.020 -34.520 1231.020 -34.510 ;
        RECT 1408.020 -34.520 1411.020 -34.510 ;
        RECT 1588.020 -34.520 1591.020 -34.510 ;
        RECT 1768.020 -34.520 1771.020 -34.510 ;
        RECT 1948.020 -34.520 1951.020 -34.510 ;
        RECT 2128.020 -34.520 2131.020 -34.510 ;
        RECT 2308.020 -34.520 2311.020 -34.510 ;
        RECT 2488.020 -34.520 2491.020 -34.510 ;
        RECT 2668.020 -34.520 2671.020 -34.510 ;
        RECT 2848.020 -34.520 2851.020 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 148.020 -37.530 151.020 -37.520 ;
        RECT 328.020 -37.530 331.020 -37.520 ;
        RECT 508.020 -37.530 511.020 -37.520 ;
        RECT 688.020 -37.530 691.020 -37.520 ;
        RECT 868.020 -37.530 871.020 -37.520 ;
        RECT 1048.020 -37.530 1051.020 -37.520 ;
        RECT 1228.020 -37.530 1231.020 -37.520 ;
        RECT 1408.020 -37.530 1411.020 -37.520 ;
        RECT 1588.020 -37.530 1591.020 -37.520 ;
        RECT 1768.020 -37.530 1771.020 -37.520 ;
        RECT 1948.020 -37.530 1951.020 -37.520 ;
        RECT 2128.020 -37.530 2131.020 -37.520 ;
        RECT 2308.020 -37.530 2311.020 -37.520 ;
        RECT 2488.020 -37.530 2491.020 -37.520 ;
        RECT 2668.020 -37.530 2671.020 -37.520 ;
        RECT 2848.020 -37.530 2851.020 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 277.840 472.555 1466.480 1449.205 ;
        RECT 1776.600 932.235 1965.200 1109.205 ;
      LAYER li1 ;
        RECT 1968.485 990.165 1968.655 1014.135 ;
      LAYER mcon ;
        RECT 1968.485 1013.965 1968.655 1014.135 ;
      LAYER met1 ;
        RECT 627.050 1473.120 627.370 1473.180 ;
        RECT 1473.450 1473.120 1473.770 1473.180 ;
        RECT 627.050 1472.980 1473.770 1473.120 ;
        RECT 627.050 1472.920 627.370 1472.980 ;
        RECT 1473.450 1472.920 1473.770 1472.980 ;
        RECT 1349.250 1472.780 1349.570 1472.840 ;
        RECT 1548.890 1472.780 1549.210 1472.840 ;
        RECT 1349.250 1472.640 1549.210 1472.780 ;
        RECT 1349.250 1472.580 1349.570 1472.640 ;
        RECT 1548.890 1472.580 1549.210 1472.640 ;
        RECT 1108.210 1472.440 1108.530 1472.500 ;
        RECT 1562.690 1472.440 1563.010 1472.500 ;
        RECT 1108.210 1472.300 1563.010 1472.440 ;
        RECT 1108.210 1472.240 1108.530 1472.300 ;
        RECT 1562.690 1472.240 1563.010 1472.300 ;
        RECT 1228.730 1472.100 1229.050 1472.160 ;
        RECT 1831.790 1472.100 1832.110 1472.160 ;
        RECT 1228.730 1471.960 1832.110 1472.100 ;
        RECT 1228.730 1471.900 1229.050 1471.960 ;
        RECT 1831.790 1471.900 1832.110 1471.960 ;
        RECT 987.690 1471.760 988.010 1471.820 ;
        RECT 1604.090 1471.760 1604.410 1471.820 ;
        RECT 987.690 1471.620 1604.410 1471.760 ;
        RECT 987.690 1471.560 988.010 1471.620 ;
        RECT 1604.090 1471.560 1604.410 1471.620 ;
        RECT 868.090 1471.420 868.410 1471.480 ;
        RECT 1610.990 1471.420 1611.310 1471.480 ;
        RECT 868.090 1471.280 1611.310 1471.420 ;
        RECT 868.090 1471.220 868.410 1471.280 ;
        RECT 1610.990 1471.220 1611.310 1471.280 ;
        RECT 747.570 1471.080 747.890 1471.140 ;
        RECT 1541.990 1471.080 1542.310 1471.140 ;
        RECT 747.570 1470.940 1542.310 1471.080 ;
        RECT 747.570 1470.880 747.890 1470.940 ;
        RECT 1541.990 1470.880 1542.310 1470.940 ;
        RECT 1468.850 1470.740 1469.170 1470.800 ;
        RECT 1968.870 1470.740 1969.190 1470.800 ;
        RECT 1468.850 1470.600 1969.190 1470.740 ;
        RECT 1468.850 1470.540 1469.170 1470.600 ;
        RECT 1968.870 1470.540 1969.190 1470.600 ;
        RECT 506.530 1470.400 506.850 1470.460 ;
        RECT 1787.170 1470.400 1787.490 1470.460 ;
        RECT 506.530 1470.260 1787.490 1470.400 ;
        RECT 506.530 1470.200 506.850 1470.260 ;
        RECT 1787.170 1470.200 1787.490 1470.260 ;
        RECT 386.930 1470.060 387.250 1470.120 ;
        RECT 1811.090 1470.060 1811.410 1470.120 ;
        RECT 386.930 1469.920 1811.410 1470.060 ;
        RECT 386.930 1469.860 387.250 1469.920 ;
        RECT 1811.090 1469.860 1811.410 1469.920 ;
        RECT 275.150 1452.040 275.470 1452.100 ;
        RECT 1980.370 1452.040 1980.690 1452.100 ;
        RECT 275.150 1451.900 1980.690 1452.040 ;
        RECT 275.150 1451.840 275.470 1451.900 ;
        RECT 1980.370 1451.840 1980.690 1451.900 ;
      LAYER met1 ;
        RECT 277.840 472.400 1468.250 1451.460 ;
      LAYER met1 ;
        RECT 1811.090 1135.840 1811.410 1135.900 ;
        RECT 1861.690 1135.840 1862.010 1135.900 ;
        RECT 1811.090 1135.700 1862.010 1135.840 ;
        RECT 1811.090 1135.640 1811.410 1135.700 ;
        RECT 1861.690 1135.640 1862.010 1135.700 ;
        RECT 1831.790 1135.160 1832.110 1135.220 ;
        RECT 1944.490 1135.160 1944.810 1135.220 ;
        RECT 1831.790 1135.020 1944.810 1135.160 ;
        RECT 1831.790 1134.960 1832.110 1135.020 ;
        RECT 1944.490 1134.960 1944.810 1135.020 ;
        RECT 1583.390 1132.100 1583.710 1132.160 ;
        RECT 1779.810 1132.100 1780.130 1132.160 ;
        RECT 1583.390 1131.960 1780.130 1132.100 ;
        RECT 1583.390 1131.900 1583.710 1131.960 ;
        RECT 1779.810 1131.900 1780.130 1131.960 ;
        RECT 1617.890 1131.760 1618.210 1131.820 ;
        RECT 1967.490 1131.760 1967.810 1131.820 ;
        RECT 1617.890 1131.620 1967.810 1131.760 ;
        RECT 1617.890 1131.560 1618.210 1131.620 ;
        RECT 1967.490 1131.560 1967.810 1131.620 ;
        RECT 1521.290 1104.220 1521.610 1104.280 ;
        RECT 1752.670 1104.220 1752.990 1104.280 ;
        RECT 1521.290 1104.080 1752.990 1104.220 ;
        RECT 1521.290 1104.020 1521.610 1104.080 ;
        RECT 1752.670 1104.020 1752.990 1104.080 ;
        RECT 1610.990 1089.940 1611.310 1090.000 ;
        RECT 1752.670 1089.940 1752.990 1090.000 ;
        RECT 1610.990 1089.800 1752.990 1089.940 ;
        RECT 1610.990 1089.740 1611.310 1089.800 ;
        RECT 1752.670 1089.740 1752.990 1089.800 ;
        RECT 1487.250 1049.140 1487.570 1049.200 ;
        RECT 1752.670 1049.140 1752.990 1049.200 ;
        RECT 1487.250 1049.000 1752.990 1049.140 ;
        RECT 1487.250 1048.940 1487.570 1049.000 ;
        RECT 1752.670 1048.940 1752.990 1049.000 ;
        RECT 1493.690 1014.460 1494.010 1014.520 ;
        RECT 1752.670 1014.460 1752.990 1014.520 ;
        RECT 1493.690 1014.320 1752.990 1014.460 ;
        RECT 1493.690 1014.260 1494.010 1014.320 ;
        RECT 1752.670 1014.260 1752.990 1014.320 ;
      LAYER met1 ;
        RECT 1776.600 932.080 1967.890 1109.360 ;
      LAYER met1 ;
        RECT 1968.410 1014.120 1968.730 1014.180 ;
        RECT 1968.215 1013.980 1968.730 1014.120 ;
        RECT 1968.410 1013.920 1968.730 1013.980 ;
        RECT 1968.410 990.320 1968.730 990.380 ;
        RECT 1968.215 990.180 1968.730 990.320 ;
        RECT 1968.410 990.120 1968.730 990.180 ;
        RECT 1487.710 931.840 1488.030 931.900 ;
        RECT 1752.670 931.840 1752.990 931.900 ;
        RECT 1487.710 931.700 1752.990 931.840 ;
        RECT 1487.710 931.640 1488.030 931.700 ;
        RECT 1752.670 931.640 1752.990 931.700 ;
        RECT 1488.170 910.760 1488.490 910.820 ;
        RECT 1956.450 910.760 1956.770 910.820 ;
        RECT 1488.170 910.620 1956.770 910.760 ;
        RECT 1488.170 910.560 1488.490 910.620 ;
        RECT 1956.450 910.560 1956.770 910.620 ;
        RECT 1548.890 910.080 1549.210 910.140 ;
        RECT 1944.490 910.080 1944.810 910.140 ;
        RECT 1548.890 909.940 1944.810 910.080 ;
        RECT 1548.890 909.880 1549.210 909.940 ;
        RECT 1944.490 909.880 1944.810 909.940 ;
        RECT 1541.990 909.740 1542.310 909.800 ;
        RECT 1921.490 909.740 1921.810 909.800 ;
        RECT 1541.990 909.600 1921.810 909.740 ;
        RECT 1541.990 909.540 1542.310 909.600 ;
        RECT 1921.490 909.540 1921.810 909.600 ;
        RECT 1486.790 909.400 1487.110 909.460 ;
        RECT 1862.610 909.400 1862.930 909.460 ;
        RECT 1486.790 909.260 1862.930 909.400 ;
        RECT 1486.790 909.200 1487.110 909.260 ;
        RECT 1862.610 909.200 1862.930 909.260 ;
        RECT 1473.450 909.060 1473.770 909.120 ;
        RECT 1776.590 909.060 1776.910 909.120 ;
        RECT 1791.770 909.060 1792.090 909.120 ;
        RECT 1473.450 908.920 1776.360 909.060 ;
        RECT 1473.450 908.860 1473.770 908.920 ;
        RECT 1776.220 908.720 1776.360 908.920 ;
        RECT 1776.590 908.920 1792.090 909.060 ;
        RECT 1776.590 908.860 1776.910 908.920 ;
        RECT 1791.770 908.860 1792.090 908.920 ;
        RECT 1803.730 908.720 1804.050 908.780 ;
        RECT 1776.220 908.580 1804.050 908.720 ;
        RECT 1803.730 908.520 1804.050 908.580 ;
        RECT 1562.690 908.380 1563.010 908.440 ;
        RECT 1873.650 908.380 1873.970 908.440 ;
        RECT 1562.690 908.240 1873.970 908.380 ;
        RECT 1562.690 908.180 1563.010 908.240 ;
        RECT 1873.650 908.180 1873.970 908.240 ;
        RECT 1604.090 908.040 1604.410 908.100 ;
        RECT 1885.610 908.040 1885.930 908.100 ;
        RECT 1604.090 907.900 1885.930 908.040 ;
        RECT 1604.090 907.840 1604.410 907.900 ;
        RECT 1885.610 907.840 1885.930 907.900 ;
        RECT 1487.250 907.360 1487.570 907.420 ;
        RECT 1838.690 907.360 1839.010 907.420 ;
        RECT 1487.250 907.220 1839.010 907.360 ;
        RECT 1487.250 907.160 1487.570 907.220 ;
        RECT 1838.690 907.160 1839.010 907.220 ;
        RECT 1811.090 907.020 1811.410 907.080 ;
        RECT 1909.530 907.020 1909.850 907.080 ;
        RECT 1811.090 906.880 1909.850 907.020 ;
        RECT 1811.090 906.820 1811.410 906.880 ;
        RECT 1909.530 906.820 1909.850 906.880 ;
        RECT 1797.290 906.680 1797.610 906.740 ;
        RECT 1850.650 906.680 1850.970 906.740 ;
        RECT 1797.290 906.540 1850.970 906.680 ;
        RECT 1797.290 906.480 1797.610 906.540 ;
        RECT 1850.650 906.480 1850.970 906.540 ;
        RECT 335.410 448.360 335.730 448.420 ;
        RECT 1968.410 448.360 1968.730 448.420 ;
        RECT 335.410 448.220 1968.730 448.360 ;
        RECT 335.410 448.160 335.730 448.220 ;
        RECT 1968.410 448.160 1968.730 448.220 ;
        RECT 575.530 448.020 575.850 448.080 ;
        RECT 1797.290 448.020 1797.610 448.080 ;
        RECT 575.530 447.880 1797.610 448.020 ;
        RECT 575.530 447.820 575.850 447.880 ;
        RECT 1797.290 447.820 1797.610 447.880 ;
        RECT 455.930 447.680 456.250 447.740 ;
        RECT 1521.290 447.680 1521.610 447.740 ;
        RECT 455.930 447.540 1521.610 447.680 ;
        RECT 455.930 447.480 456.250 447.540 ;
        RECT 1521.290 447.480 1521.610 447.540 ;
        RECT 816.570 447.340 816.890 447.400 ;
        RECT 1776.590 447.340 1776.910 447.400 ;
        RECT 816.570 447.200 1776.910 447.340 ;
        RECT 816.570 447.140 816.890 447.200 ;
        RECT 1776.590 447.140 1776.910 447.200 ;
        RECT 696.050 447.000 696.370 447.060 ;
        RECT 1583.390 447.000 1583.710 447.060 ;
        RECT 696.050 446.860 1583.710 447.000 ;
        RECT 696.050 446.800 696.370 446.860 ;
        RECT 1583.390 446.800 1583.710 446.860 ;
        RECT 1177.210 446.660 1177.530 446.720 ;
        RECT 1969.330 446.660 1969.650 446.720 ;
        RECT 1177.210 446.520 1969.650 446.660 ;
        RECT 1177.210 446.460 1177.530 446.520 ;
        RECT 1969.330 446.460 1969.650 446.520 ;
        RECT 937.090 446.320 937.410 446.380 ;
        RECT 1617.890 446.320 1618.210 446.380 ;
        RECT 937.090 446.180 1618.210 446.320 ;
        RECT 937.090 446.120 937.410 446.180 ;
        RECT 1617.890 446.120 1618.210 446.180 ;
        RECT 1297.730 445.980 1298.050 446.040 ;
        RECT 1967.950 445.980 1968.270 446.040 ;
        RECT 1297.730 445.840 1968.270 445.980 ;
        RECT 1297.730 445.780 1298.050 445.840 ;
        RECT 1967.950 445.780 1968.270 445.840 ;
        RECT 1057.610 445.640 1057.930 445.700 ;
        RECT 1493.690 445.640 1494.010 445.700 ;
        RECT 1057.610 445.500 1494.010 445.640 ;
        RECT 1057.610 445.440 1057.930 445.500 ;
        RECT 1493.690 445.440 1494.010 445.500 ;
        RECT 1418.250 445.300 1418.570 445.360 ;
        RECT 1811.090 445.300 1811.410 445.360 ;
        RECT 1418.250 445.160 1811.410 445.300 ;
        RECT 1418.250 445.100 1418.570 445.160 ;
        RECT 1811.090 445.100 1811.410 445.160 ;
      LAYER via ;
        RECT 627.080 1472.920 627.340 1473.180 ;
        RECT 1473.480 1472.920 1473.740 1473.180 ;
        RECT 1349.280 1472.580 1349.540 1472.840 ;
        RECT 1548.920 1472.580 1549.180 1472.840 ;
        RECT 1108.240 1472.240 1108.500 1472.500 ;
        RECT 1562.720 1472.240 1562.980 1472.500 ;
        RECT 1228.760 1471.900 1229.020 1472.160 ;
        RECT 1831.820 1471.900 1832.080 1472.160 ;
        RECT 987.720 1471.560 987.980 1471.820 ;
        RECT 1604.120 1471.560 1604.380 1471.820 ;
        RECT 868.120 1471.220 868.380 1471.480 ;
        RECT 1611.020 1471.220 1611.280 1471.480 ;
        RECT 747.600 1470.880 747.860 1471.140 ;
        RECT 1542.020 1470.880 1542.280 1471.140 ;
        RECT 1468.880 1470.540 1469.140 1470.800 ;
        RECT 1968.900 1470.540 1969.160 1470.800 ;
        RECT 506.560 1470.200 506.820 1470.460 ;
        RECT 1787.200 1470.200 1787.460 1470.460 ;
        RECT 386.960 1469.860 387.220 1470.120 ;
        RECT 1811.120 1469.860 1811.380 1470.120 ;
        RECT 275.180 1451.840 275.440 1452.100 ;
        RECT 1980.400 1451.840 1980.660 1452.100 ;
        RECT 1811.120 1135.640 1811.380 1135.900 ;
        RECT 1861.720 1135.640 1861.980 1135.900 ;
        RECT 1831.820 1134.960 1832.080 1135.220 ;
        RECT 1944.520 1134.960 1944.780 1135.220 ;
        RECT 1583.420 1131.900 1583.680 1132.160 ;
        RECT 1779.840 1131.900 1780.100 1132.160 ;
        RECT 1617.920 1131.560 1618.180 1131.820 ;
        RECT 1967.520 1131.560 1967.780 1131.820 ;
        RECT 1521.320 1104.020 1521.580 1104.280 ;
        RECT 1752.700 1104.020 1752.960 1104.280 ;
        RECT 1611.020 1089.740 1611.280 1090.000 ;
        RECT 1752.700 1089.740 1752.960 1090.000 ;
        RECT 1487.280 1048.940 1487.540 1049.200 ;
        RECT 1752.700 1048.940 1752.960 1049.200 ;
        RECT 1493.720 1014.260 1493.980 1014.520 ;
        RECT 1752.700 1014.260 1752.960 1014.520 ;
        RECT 1968.440 1013.920 1968.700 1014.180 ;
        RECT 1968.440 990.120 1968.700 990.380 ;
        RECT 1487.740 931.640 1488.000 931.900 ;
        RECT 1752.700 931.640 1752.960 931.900 ;
        RECT 1488.200 910.560 1488.460 910.820 ;
        RECT 1956.480 910.560 1956.740 910.820 ;
        RECT 1548.920 909.880 1549.180 910.140 ;
        RECT 1944.520 909.880 1944.780 910.140 ;
        RECT 1542.020 909.540 1542.280 909.800 ;
        RECT 1921.520 909.540 1921.780 909.800 ;
        RECT 1486.820 909.200 1487.080 909.460 ;
        RECT 1862.640 909.200 1862.900 909.460 ;
        RECT 1473.480 908.860 1473.740 909.120 ;
        RECT 1776.620 908.860 1776.880 909.120 ;
        RECT 1791.800 908.860 1792.060 909.120 ;
        RECT 1803.760 908.520 1804.020 908.780 ;
        RECT 1562.720 908.180 1562.980 908.440 ;
        RECT 1873.680 908.180 1873.940 908.440 ;
        RECT 1604.120 907.840 1604.380 908.100 ;
        RECT 1885.640 907.840 1885.900 908.100 ;
        RECT 1487.280 907.160 1487.540 907.420 ;
        RECT 1838.720 907.160 1838.980 907.420 ;
        RECT 1811.120 906.820 1811.380 907.080 ;
        RECT 1909.560 906.820 1909.820 907.080 ;
        RECT 1797.320 906.480 1797.580 906.740 ;
        RECT 1850.680 906.480 1850.940 906.740 ;
        RECT 335.440 448.160 335.700 448.420 ;
        RECT 1968.440 448.160 1968.700 448.420 ;
        RECT 575.560 447.820 575.820 448.080 ;
        RECT 1797.320 447.820 1797.580 448.080 ;
        RECT 455.960 447.480 456.220 447.740 ;
        RECT 1521.320 447.480 1521.580 447.740 ;
        RECT 816.600 447.140 816.860 447.400 ;
        RECT 1776.620 447.140 1776.880 447.400 ;
        RECT 696.080 446.800 696.340 447.060 ;
        RECT 1583.420 446.800 1583.680 447.060 ;
        RECT 1177.240 446.460 1177.500 446.720 ;
        RECT 1969.360 446.460 1969.620 446.720 ;
        RECT 937.120 446.120 937.380 446.380 ;
        RECT 1617.920 446.120 1618.180 446.380 ;
        RECT 1297.760 445.780 1298.020 446.040 ;
        RECT 1967.980 445.780 1968.240 446.040 ;
        RECT 1057.640 445.440 1057.900 445.700 ;
        RECT 1493.720 445.440 1493.980 445.700 ;
        RECT 1418.280 445.100 1418.540 445.360 ;
        RECT 1811.120 445.100 1811.380 445.360 ;
      LAYER met2 ;
        RECT 627.080 1472.890 627.340 1473.210 ;
        RECT 1473.480 1472.890 1473.740 1473.210 ;
        RECT 506.560 1470.170 506.820 1470.490 ;
        RECT 386.960 1469.830 387.220 1470.150 ;
        RECT 387.020 1460.000 387.160 1469.830 ;
        RECT 506.620 1460.000 506.760 1470.170 ;
        RECT 627.140 1460.000 627.280 1472.890 ;
        RECT 1349.280 1472.550 1349.540 1472.870 ;
        RECT 1108.240 1472.210 1108.500 1472.530 ;
        RECT 987.720 1471.530 987.980 1471.850 ;
        RECT 868.120 1471.190 868.380 1471.510 ;
        RECT 747.600 1470.850 747.860 1471.170 ;
        RECT 747.660 1460.000 747.800 1470.850 ;
        RECT 868.180 1460.000 868.320 1471.190 ;
        RECT 987.780 1460.000 987.920 1471.530 ;
        RECT 1108.300 1460.000 1108.440 1472.210 ;
        RECT 1228.760 1471.870 1229.020 1472.190 ;
        RECT 1228.820 1460.000 1228.960 1471.870 ;
        RECT 1349.340 1460.000 1349.480 1472.550 ;
        RECT 1468.880 1470.510 1469.140 1470.830 ;
        RECT 1468.940 1460.000 1469.080 1470.510 ;
        RECT 386.950 1456.000 387.230 1460.000 ;
        RECT 506.550 1456.000 506.830 1460.000 ;
        RECT 627.070 1456.000 627.350 1460.000 ;
        RECT 747.590 1456.000 747.870 1460.000 ;
        RECT 868.110 1456.000 868.390 1460.000 ;
        RECT 987.710 1456.000 987.990 1460.000 ;
        RECT 1108.230 1456.000 1108.510 1460.000 ;
        RECT 1228.750 1456.000 1229.030 1460.000 ;
        RECT 1349.270 1456.000 1349.550 1460.000 ;
        RECT 1468.870 1456.000 1469.150 1460.000 ;
      LAYER met2 ;
        RECT 280.700 1455.720 386.670 1456.000 ;
        RECT 387.510 1455.720 506.270 1456.000 ;
        RECT 507.110 1455.720 626.790 1456.000 ;
        RECT 627.630 1455.720 747.310 1456.000 ;
        RECT 748.150 1455.720 867.830 1456.000 ;
        RECT 868.670 1455.720 987.430 1456.000 ;
        RECT 988.270 1455.720 1107.950 1456.000 ;
        RECT 1108.790 1455.720 1228.470 1456.000 ;
        RECT 1229.310 1455.720 1348.990 1456.000 ;
        RECT 1349.830 1455.720 1468.590 1456.000 ;
        RECT 1469.430 1455.720 1470.070 1456.000 ;
      LAYER met2 ;
        RECT 275.180 1451.810 275.440 1452.130 ;
        RECT 275.240 1446.205 275.380 1451.810 ;
        RECT 275.170 1445.835 275.450 1446.205 ;
        RECT 261.830 553.675 262.110 554.045 ;
        RECT 261.900 471.765 262.040 553.675 ;
        RECT 261.830 471.395 262.110 471.765 ;
      LAYER met2 ;
        RECT 280.700 464.280 1470.070 1455.720 ;
      LAYER met2 ;
        RECT 1473.540 909.150 1473.680 1472.890 ;
        RECT 1548.920 1472.550 1549.180 1472.870 ;
        RECT 1542.020 1470.850 1542.280 1471.170 ;
        RECT 1486.810 1278.555 1487.090 1278.925 ;
        RECT 1486.880 909.490 1487.020 1278.555 ;
        RECT 1521.320 1103.990 1521.580 1104.310 ;
        RECT 1488.190 1100.395 1488.470 1100.765 ;
        RECT 1487.280 1048.910 1487.540 1049.230 ;
        RECT 1487.340 922.605 1487.480 1048.910 ;
        RECT 1487.740 931.610 1488.000 931.930 ;
        RECT 1487.270 922.235 1487.550 922.605 ;
        RECT 1486.820 909.170 1487.080 909.490 ;
        RECT 1473.480 908.830 1473.740 909.150 ;
        RECT 1487.280 907.130 1487.540 907.450 ;
        RECT 1487.340 567.645 1487.480 907.130 ;
        RECT 1487.800 744.445 1487.940 931.610 ;
        RECT 1488.260 910.850 1488.400 1100.395 ;
        RECT 1493.720 1014.230 1493.980 1014.550 ;
        RECT 1488.200 910.530 1488.460 910.850 ;
        RECT 1487.730 744.075 1488.010 744.445 ;
        RECT 1487.270 567.275 1487.550 567.645 ;
      LAYER met2 ;
        RECT 280.700 464.000 335.150 464.280 ;
        RECT 335.990 464.000 455.670 464.280 ;
        RECT 456.510 464.000 575.270 464.280 ;
        RECT 576.110 464.000 695.790 464.280 ;
        RECT 696.630 464.000 816.310 464.280 ;
        RECT 817.150 464.000 936.830 464.280 ;
        RECT 937.670 464.000 1057.350 464.280 ;
        RECT 1058.190 464.000 1176.950 464.280 ;
        RECT 1177.790 464.000 1297.470 464.280 ;
        RECT 1298.310 464.000 1417.990 464.280 ;
        RECT 1418.830 464.000 1470.070 464.280 ;
      LAYER met2 ;
        RECT 335.430 460.000 335.710 464.000 ;
        RECT 455.950 460.000 456.230 464.000 ;
        RECT 575.550 460.000 575.830 464.000 ;
        RECT 696.070 460.000 696.350 464.000 ;
        RECT 816.590 460.000 816.870 464.000 ;
        RECT 937.110 460.000 937.390 464.000 ;
        RECT 1057.630 460.000 1057.910 464.000 ;
        RECT 1177.230 460.000 1177.510 464.000 ;
        RECT 1297.750 460.000 1298.030 464.000 ;
        RECT 1418.270 460.000 1418.550 464.000 ;
        RECT 335.500 448.450 335.640 460.000 ;
        RECT 335.440 448.130 335.700 448.450 ;
        RECT 456.020 447.770 456.160 460.000 ;
        RECT 575.620 448.110 575.760 460.000 ;
        RECT 575.560 447.790 575.820 448.110 ;
        RECT 455.960 447.450 456.220 447.770 ;
        RECT 696.140 447.090 696.280 460.000 ;
        RECT 816.660 447.430 816.800 460.000 ;
        RECT 816.600 447.110 816.860 447.430 ;
        RECT 696.080 446.770 696.340 447.090 ;
        RECT 937.180 446.410 937.320 460.000 ;
        RECT 937.120 446.090 937.380 446.410 ;
        RECT 1057.700 445.730 1057.840 460.000 ;
        RECT 1177.300 446.750 1177.440 460.000 ;
        RECT 1177.240 446.430 1177.500 446.750 ;
        RECT 1297.820 446.070 1297.960 460.000 ;
        RECT 1297.760 445.750 1298.020 446.070 ;
        RECT 1057.640 445.410 1057.900 445.730 ;
        RECT 1418.340 445.390 1418.480 460.000 ;
        RECT 1493.780 445.730 1493.920 1014.230 ;
        RECT 1521.380 447.770 1521.520 1103.990 ;
        RECT 1542.080 909.830 1542.220 1470.850 ;
        RECT 1548.980 910.170 1549.120 1472.550 ;
        RECT 1562.720 1472.210 1562.980 1472.530 ;
        RECT 1548.920 909.850 1549.180 910.170 ;
        RECT 1542.020 909.510 1542.280 909.830 ;
        RECT 1562.780 908.470 1562.920 1472.210 ;
        RECT 1831.820 1471.870 1832.080 1472.190 ;
        RECT 1604.120 1471.530 1604.380 1471.850 ;
        RECT 1583.420 1131.870 1583.680 1132.190 ;
        RECT 1562.720 908.150 1562.980 908.470 ;
        RECT 1521.320 447.450 1521.580 447.770 ;
        RECT 1583.480 447.090 1583.620 1131.870 ;
        RECT 1604.180 908.130 1604.320 1471.530 ;
        RECT 1611.020 1471.190 1611.280 1471.510 ;
        RECT 1611.080 1090.030 1611.220 1471.190 ;
        RECT 1787.200 1470.170 1787.460 1470.490 ;
        RECT 1779.840 1131.870 1780.100 1132.190 ;
        RECT 1617.920 1131.530 1618.180 1131.850 ;
        RECT 1611.020 1089.710 1611.280 1090.030 ;
        RECT 1604.120 907.810 1604.380 908.130 ;
        RECT 1583.420 446.770 1583.680 447.090 ;
        RECT 1617.980 446.410 1618.120 1131.530 ;
        RECT 1779.900 1120.000 1780.040 1131.870 ;
        RECT 1787.260 1120.370 1787.400 1470.170 ;
        RECT 1811.120 1469.830 1811.380 1470.150 ;
        RECT 1811.180 1135.930 1811.320 1469.830 ;
        RECT 1811.120 1135.610 1811.380 1135.930 ;
        RECT 1831.880 1135.250 1832.020 1471.870 ;
        RECT 1968.900 1470.510 1969.160 1470.830 ;
        RECT 1861.720 1135.610 1861.980 1135.930 ;
        RECT 1831.820 1134.930 1832.080 1135.250 ;
        RECT 1838.710 1133.715 1838.990 1134.085 ;
        RECT 1826.750 1131.675 1827.030 1132.045 ;
        RECT 1787.260 1120.230 1789.700 1120.370 ;
        RECT 1779.900 1119.620 1780.190 1120.000 ;
        RECT 1779.910 1116.000 1780.190 1119.620 ;
        RECT 1789.560 1119.690 1789.700 1120.230 ;
        RECT 1826.820 1120.000 1826.960 1131.675 ;
        RECT 1838.780 1120.000 1838.920 1133.715 ;
        RECT 1861.780 1120.000 1861.920 1135.610 ;
        RECT 1944.520 1134.930 1944.780 1135.250 ;
        RECT 1944.580 1120.000 1944.720 1134.930 ;
        RECT 1967.520 1131.530 1967.780 1131.850 ;
        RECT 1967.580 1120.000 1967.720 1131.530 ;
        RECT 1790.950 1119.690 1791.230 1120.000 ;
        RECT 1789.560 1119.550 1791.230 1119.690 ;
        RECT 1826.820 1119.620 1827.110 1120.000 ;
        RECT 1838.780 1119.620 1839.070 1120.000 ;
        RECT 1861.780 1119.620 1862.070 1120.000 ;
        RECT 1790.950 1116.000 1791.230 1119.550 ;
        RECT 1826.830 1116.000 1827.110 1119.620 ;
        RECT 1838.790 1116.000 1839.070 1119.620 ;
        RECT 1861.790 1116.000 1862.070 1119.620 ;
        RECT 1907.250 1118.330 1907.530 1118.445 ;
        RECT 1908.710 1118.330 1908.990 1120.000 ;
        RECT 1907.250 1118.190 1908.990 1118.330 ;
        RECT 1907.250 1118.075 1907.530 1118.190 ;
        RECT 1908.710 1116.000 1908.990 1118.190 ;
        RECT 1919.210 1118.330 1919.490 1118.445 ;
        RECT 1920.670 1118.330 1920.950 1120.000 ;
        RECT 1944.580 1119.620 1944.870 1120.000 ;
        RECT 1967.580 1119.620 1967.870 1120.000 ;
        RECT 1919.210 1118.190 1920.950 1118.330 ;
        RECT 1919.210 1118.075 1919.490 1118.190 ;
        RECT 1920.670 1116.000 1920.950 1118.190 ;
        RECT 1944.590 1116.000 1944.870 1119.620 ;
        RECT 1967.590 1116.000 1967.870 1119.620 ;
      LAYER met2 ;
        RECT 1780.470 1115.720 1790.670 1116.000 ;
        RECT 1791.510 1115.720 1802.630 1116.000 ;
        RECT 1803.470 1115.720 1814.590 1116.000 ;
        RECT 1815.430 1115.720 1826.550 1116.000 ;
        RECT 1827.390 1115.720 1838.510 1116.000 ;
        RECT 1839.350 1115.720 1849.550 1116.000 ;
        RECT 1850.390 1115.720 1861.510 1116.000 ;
        RECT 1862.350 1115.720 1873.470 1116.000 ;
        RECT 1874.310 1115.720 1885.430 1116.000 ;
        RECT 1886.270 1115.720 1897.390 1116.000 ;
        RECT 1898.230 1115.720 1908.430 1116.000 ;
        RECT 1909.270 1115.720 1920.390 1116.000 ;
        RECT 1921.230 1115.720 1932.350 1116.000 ;
        RECT 1933.190 1115.720 1944.310 1116.000 ;
        RECT 1945.150 1115.720 1956.270 1116.000 ;
        RECT 1957.110 1115.720 1967.310 1116.000 ;
      LAYER met2 ;
        RECT 1752.690 1107.195 1752.970 1107.565 ;
        RECT 1752.760 1104.310 1752.900 1107.195 ;
        RECT 1752.700 1103.990 1752.960 1104.310 ;
        RECT 1752.700 1089.885 1752.960 1090.030 ;
        RECT 1752.690 1089.515 1752.970 1089.885 ;
        RECT 1752.690 1054.155 1752.970 1054.525 ;
        RECT 1752.760 1049.230 1752.900 1054.155 ;
        RECT 1752.700 1048.910 1752.960 1049.230 ;
        RECT 1752.690 1020.155 1752.970 1020.525 ;
        RECT 1752.760 1014.550 1752.900 1020.155 ;
        RECT 1752.700 1014.230 1752.960 1014.550 ;
        RECT 1752.690 933.115 1752.970 933.485 ;
        RECT 1752.760 931.930 1752.900 933.115 ;
        RECT 1752.700 931.610 1752.960 931.930 ;
      LAYER met2 ;
        RECT 1779.920 924.280 1967.860 1115.720 ;
      LAYER met2 ;
        RECT 1968.430 1078.635 1968.710 1079.005 ;
        RECT 1968.500 1014.210 1968.640 1078.635 ;
        RECT 1968.960 1014.970 1969.100 1470.510 ;
        RECT 1980.400 1451.810 1980.660 1452.130 ;
        RECT 1980.460 1099.405 1980.600 1451.810 ;
        RECT 1980.390 1099.035 1980.670 1099.405 ;
        RECT 1968.960 1014.830 1970.480 1014.970 ;
        RECT 1968.440 1013.890 1968.700 1014.210 ;
        RECT 1968.430 993.210 1968.710 993.325 ;
      LAYER met2 ;
        RECT 1780.470 924.000 1791.590 924.280 ;
        RECT 1792.430 924.000 1803.550 924.280 ;
        RECT 1804.390 924.000 1814.590 924.280 ;
        RECT 1815.430 924.000 1826.550 924.280 ;
        RECT 1827.390 924.000 1838.510 924.280 ;
        RECT 1839.350 924.000 1850.470 924.280 ;
        RECT 1851.310 924.000 1862.430 924.280 ;
        RECT 1863.270 924.000 1873.470 924.280 ;
        RECT 1874.310 924.000 1885.430 924.280 ;
        RECT 1886.270 924.000 1897.390 924.280 ;
        RECT 1898.230 924.000 1909.350 924.280 ;
        RECT 1910.190 924.000 1921.310 924.280 ;
        RECT 1922.150 924.000 1932.350 924.280 ;
        RECT 1933.190 924.000 1944.310 924.280 ;
        RECT 1945.150 924.000 1956.270 924.280 ;
        RECT 1957.110 924.000 1967.860 924.280 ;
      LAYER met2 ;
        RECT 1968.040 993.070 1968.710 993.210 ;
        RECT 1791.870 920.380 1792.150 924.000 ;
        RECT 1803.830 920.380 1804.110 924.000 ;
        RECT 1838.790 920.380 1839.070 924.000 ;
        RECT 1850.750 920.380 1851.030 924.000 ;
        RECT 1862.710 920.380 1862.990 924.000 ;
        RECT 1873.750 920.380 1874.030 924.000 ;
        RECT 1885.710 920.380 1885.990 924.000 ;
        RECT 1909.630 920.380 1909.910 924.000 ;
        RECT 1921.590 920.380 1921.870 924.000 ;
        RECT 1944.590 920.380 1944.870 924.000 ;
        RECT 1956.550 920.380 1956.830 924.000 ;
        RECT 1791.860 920.000 1792.150 920.380 ;
        RECT 1803.820 920.000 1804.110 920.380 ;
        RECT 1838.780 920.000 1839.070 920.380 ;
        RECT 1850.740 920.000 1851.030 920.380 ;
        RECT 1862.700 920.000 1862.990 920.380 ;
        RECT 1873.740 920.000 1874.030 920.380 ;
        RECT 1885.700 920.000 1885.990 920.380 ;
        RECT 1909.620 920.000 1909.910 920.380 ;
        RECT 1921.580 920.000 1921.870 920.380 ;
        RECT 1944.580 920.000 1944.870 920.380 ;
        RECT 1956.540 920.000 1956.830 920.380 ;
        RECT 1791.860 909.150 1792.000 920.000 ;
        RECT 1776.620 908.830 1776.880 909.150 ;
        RECT 1791.800 908.830 1792.060 909.150 ;
        RECT 1776.680 447.430 1776.820 908.830 ;
        RECT 1803.820 908.810 1803.960 920.000 ;
        RECT 1803.760 908.490 1804.020 908.810 ;
        RECT 1838.780 907.450 1838.920 920.000 ;
        RECT 1838.720 907.130 1838.980 907.450 ;
        RECT 1811.120 906.790 1811.380 907.110 ;
        RECT 1797.320 906.450 1797.580 906.770 ;
        RECT 1797.380 448.110 1797.520 906.450 ;
        RECT 1797.320 447.790 1797.580 448.110 ;
        RECT 1776.620 447.110 1776.880 447.430 ;
        RECT 1617.920 446.090 1618.180 446.410 ;
        RECT 1493.720 445.410 1493.980 445.730 ;
        RECT 1811.180 445.390 1811.320 906.790 ;
        RECT 1850.740 906.770 1850.880 920.000 ;
        RECT 1862.700 909.490 1862.840 920.000 ;
        RECT 1862.640 909.170 1862.900 909.490 ;
        RECT 1873.740 908.470 1873.880 920.000 ;
        RECT 1873.680 908.150 1873.940 908.470 ;
        RECT 1885.700 908.130 1885.840 920.000 ;
        RECT 1885.640 907.810 1885.900 908.130 ;
        RECT 1909.620 907.110 1909.760 920.000 ;
        RECT 1921.580 909.830 1921.720 920.000 ;
        RECT 1944.580 910.170 1944.720 920.000 ;
        RECT 1956.540 910.850 1956.680 920.000 ;
        RECT 1956.480 910.530 1956.740 910.850 ;
        RECT 1944.520 909.850 1944.780 910.170 ;
        RECT 1921.520 909.510 1921.780 909.830 ;
        RECT 1909.560 906.790 1909.820 907.110 ;
        RECT 1850.680 906.450 1850.940 906.770 ;
        RECT 1968.040 446.070 1968.180 993.070 ;
        RECT 1968.430 992.955 1968.710 993.070 ;
        RECT 1968.440 990.090 1968.700 990.410 ;
        RECT 1968.500 448.450 1968.640 990.090 ;
        RECT 1970.340 979.610 1970.480 1014.830 ;
        RECT 1968.960 979.470 1970.480 979.610 ;
        RECT 1968.960 945.045 1969.100 979.470 ;
        RECT 1969.350 973.915 1969.630 974.285 ;
        RECT 1968.890 944.675 1969.170 945.045 ;
        RECT 1968.440 448.130 1968.700 448.450 ;
        RECT 1969.420 446.750 1969.560 973.915 ;
        RECT 1969.360 446.430 1969.620 446.750 ;
        RECT 1967.980 445.750 1968.240 446.070 ;
        RECT 1418.280 445.070 1418.540 445.390 ;
        RECT 1811.120 445.070 1811.380 445.390 ;
      LAYER via2 ;
        RECT 275.170 1445.880 275.450 1446.160 ;
        RECT 261.830 553.720 262.110 554.000 ;
        RECT 261.830 471.440 262.110 471.720 ;
        RECT 1486.810 1278.600 1487.090 1278.880 ;
        RECT 1488.190 1100.440 1488.470 1100.720 ;
        RECT 1487.270 922.280 1487.550 922.560 ;
        RECT 1487.730 744.120 1488.010 744.400 ;
        RECT 1487.270 567.320 1487.550 567.600 ;
        RECT 1838.710 1133.760 1838.990 1134.040 ;
        RECT 1826.750 1131.720 1827.030 1132.000 ;
        RECT 1907.250 1118.120 1907.530 1118.400 ;
        RECT 1919.210 1118.120 1919.490 1118.400 ;
        RECT 1752.690 1107.240 1752.970 1107.520 ;
        RECT 1752.690 1089.560 1752.970 1089.840 ;
        RECT 1752.690 1054.200 1752.970 1054.480 ;
        RECT 1752.690 1020.200 1752.970 1020.480 ;
        RECT 1752.690 933.160 1752.970 933.440 ;
        RECT 1968.430 1078.680 1968.710 1078.960 ;
        RECT 1980.390 1099.080 1980.670 1099.360 ;
        RECT 1968.430 993.000 1968.710 993.280 ;
        RECT 1969.350 973.960 1969.630 974.240 ;
        RECT 1968.890 944.720 1969.170 945.000 ;
      LAYER met3 ;
        RECT 275.145 1446.170 275.475 1446.185 ;
        RECT 275.145 1445.855 275.690 1446.170 ;
        RECT 275.390 1443.640 275.690 1445.855 ;
      LAYER met3 ;
        RECT 276.000 1444.040 1471.730 1449.285 ;
      LAYER met3 ;
        RECT 272.000 1443.040 276.000 1443.640 ;
      LAYER met3 ;
        RECT 276.400 1442.640 1471.730 1444.040 ;
        RECT 276.000 1279.480 1471.730 1442.640 ;
        RECT 276.000 1278.080 1467.600 1279.480 ;
      LAYER met3 ;
        RECT 1468.000 1278.890 1472.000 1279.080 ;
        RECT 1486.785 1278.890 1487.115 1278.905 ;
        RECT 1468.000 1278.590 1487.115 1278.890 ;
        RECT 1468.000 1278.480 1472.000 1278.590 ;
        RECT 1486.785 1278.575 1487.115 1278.590 ;
      LAYER met3 ;
        RECT 276.000 1265.880 1471.730 1278.080 ;
      LAYER met3 ;
        RECT 261.550 1265.290 261.930 1265.300 ;
        RECT 272.000 1265.290 276.000 1265.480 ;
        RECT 261.550 1264.990 276.000 1265.290 ;
        RECT 261.550 1264.980 261.930 1264.990 ;
        RECT 272.000 1264.880 276.000 1264.990 ;
      LAYER met3 ;
        RECT 276.400 1264.480 1471.730 1265.880 ;
        RECT 276.000 1101.320 1471.730 1264.480 ;
      LAYER met3 ;
        RECT 1545.870 1140.850 1546.250 1140.860 ;
        RECT 1592.790 1140.850 1593.170 1140.860 ;
        RECT 1545.870 1140.550 1593.170 1140.850 ;
        RECT 1545.870 1140.540 1546.250 1140.550 ;
        RECT 1592.790 1140.540 1593.170 1140.550 ;
        RECT 1646.150 1140.850 1646.530 1140.860 ;
        RECT 1689.390 1140.850 1689.770 1140.860 ;
        RECT 1646.150 1140.550 1689.770 1140.850 ;
        RECT 1646.150 1140.540 1646.530 1140.550 ;
        RECT 1689.390 1140.540 1689.770 1140.550 ;
        RECT 1739.070 1140.850 1739.450 1140.860 ;
        RECT 1785.990 1140.850 1786.370 1140.860 ;
        RECT 1739.070 1140.550 1786.370 1140.850 ;
        RECT 1739.070 1140.540 1739.450 1140.550 ;
        RECT 1785.990 1140.540 1786.370 1140.550 ;
        RECT 1800.710 1134.050 1801.090 1134.060 ;
        RECT 1838.685 1134.050 1839.015 1134.065 ;
        RECT 1800.710 1133.750 1839.015 1134.050 ;
        RECT 1800.710 1133.740 1801.090 1133.750 ;
        RECT 1838.685 1133.735 1839.015 1133.750 ;
        RECT 1783.230 1132.010 1783.610 1132.020 ;
        RECT 1826.725 1132.010 1827.055 1132.025 ;
        RECT 1783.230 1131.710 1827.055 1132.010 ;
        RECT 1783.230 1131.700 1783.610 1131.710 ;
        RECT 1826.725 1131.695 1827.055 1131.710 ;
        RECT 1904.670 1118.410 1905.050 1118.420 ;
        RECT 1907.225 1118.410 1907.555 1118.425 ;
        RECT 1904.670 1118.110 1907.555 1118.410 ;
        RECT 1904.670 1118.100 1905.050 1118.110 ;
        RECT 1907.225 1118.095 1907.555 1118.110 ;
        RECT 1918.470 1118.410 1918.850 1118.420 ;
        RECT 1919.185 1118.410 1919.515 1118.425 ;
        RECT 1918.470 1118.110 1919.515 1118.410 ;
        RECT 1918.470 1118.100 1918.850 1118.110 ;
        RECT 1919.185 1118.095 1919.515 1118.110 ;
      LAYER met3 ;
        RECT 1774.720 1108.120 1966.720 1109.285 ;
      LAYER met3 ;
        RECT 1752.665 1107.530 1752.995 1107.545 ;
        RECT 1770.720 1107.530 1774.720 1107.720 ;
        RECT 1752.665 1107.230 1774.720 1107.530 ;
        RECT 1752.665 1107.215 1752.995 1107.230 ;
        RECT 1770.720 1107.120 1774.720 1107.230 ;
      LAYER met3 ;
        RECT 1775.120 1106.720 1966.720 1108.120 ;
        RECT 276.000 1099.920 1467.600 1101.320 ;
      LAYER met3 ;
        RECT 1468.000 1100.730 1472.000 1100.920 ;
        RECT 1488.165 1100.730 1488.495 1100.745 ;
        RECT 1468.000 1100.430 1488.495 1100.730 ;
        RECT 1468.000 1100.320 1472.000 1100.430 ;
        RECT 1488.165 1100.415 1488.495 1100.430 ;
      LAYER met3 ;
        RECT 1774.720 1099.960 1966.720 1106.720 ;
        RECT 276.000 1087.720 1471.730 1099.920 ;
        RECT 1774.720 1098.560 1966.320 1099.960 ;
      LAYER met3 ;
        RECT 1966.720 1099.370 1970.720 1099.560 ;
        RECT 1980.365 1099.370 1980.695 1099.385 ;
        RECT 1966.720 1099.070 1980.695 1099.370 ;
        RECT 1966.720 1098.960 1970.720 1099.070 ;
        RECT 1980.365 1099.055 1980.695 1099.070 ;
      LAYER met3 ;
        RECT 1774.720 1090.440 1966.720 1098.560 ;
      LAYER met3 ;
        RECT 1752.665 1089.850 1752.995 1089.865 ;
        RECT 1770.720 1089.850 1774.720 1090.040 ;
        RECT 1752.665 1089.550 1774.720 1089.850 ;
        RECT 1752.665 1089.535 1752.995 1089.550 ;
        RECT 1770.720 1089.440 1774.720 1089.550 ;
      LAYER met3 ;
        RECT 1775.120 1089.040 1966.720 1090.440 ;
      LAYER met3 ;
        RECT 272.000 1086.720 276.000 1087.320 ;
        RECT 272.630 1084.420 272.930 1086.720 ;
      LAYER met3 ;
        RECT 276.400 1086.320 1471.730 1087.720 ;
      LAYER met3 ;
        RECT 272.590 1084.100 272.970 1084.420 ;
      LAYER met3 ;
        RECT 276.000 923.160 1471.730 1086.320 ;
        RECT 1774.720 1082.280 1966.720 1089.040 ;
        RECT 1774.720 1080.880 1966.320 1082.280 ;
      LAYER met3 ;
        RECT 1966.720 1081.280 1970.720 1081.880 ;
      LAYER met3 ;
        RECT 1774.720 1072.760 1966.720 1080.880 ;
      LAYER met3 ;
        RECT 1968.190 1078.985 1968.490 1081.280 ;
        RECT 1968.190 1078.670 1968.735 1078.985 ;
        RECT 1968.405 1078.655 1968.735 1078.670 ;
      LAYER met3 ;
        RECT 1775.120 1071.360 1966.720 1072.760 ;
        RECT 1774.720 1064.600 1966.720 1071.360 ;
        RECT 1774.720 1063.200 1966.320 1064.600 ;
        RECT 1774.720 1055.080 1966.720 1063.200 ;
      LAYER met3 ;
        RECT 1752.665 1054.490 1752.995 1054.505 ;
        RECT 1770.720 1054.490 1774.720 1054.680 ;
        RECT 1752.665 1054.190 1774.720 1054.490 ;
        RECT 1752.665 1054.175 1752.995 1054.190 ;
        RECT 1770.720 1054.080 1774.720 1054.190 ;
      LAYER met3 ;
        RECT 1775.120 1053.680 1966.720 1055.080 ;
        RECT 1774.720 1046.920 1966.720 1053.680 ;
        RECT 1774.720 1045.520 1966.320 1046.920 ;
        RECT 1774.720 1038.760 1966.720 1045.520 ;
        RECT 1775.120 1037.360 1966.720 1038.760 ;
        RECT 1774.720 1030.600 1966.720 1037.360 ;
        RECT 1774.720 1029.200 1966.320 1030.600 ;
        RECT 1774.720 1021.080 1966.720 1029.200 ;
      LAYER met3 ;
        RECT 1752.665 1020.490 1752.995 1020.505 ;
        RECT 1770.720 1020.490 1774.720 1020.680 ;
        RECT 1752.665 1020.190 1774.720 1020.490 ;
        RECT 1752.665 1020.175 1752.995 1020.190 ;
        RECT 1770.720 1020.080 1774.720 1020.190 ;
      LAYER met3 ;
        RECT 1775.120 1019.680 1966.720 1021.080 ;
        RECT 1774.720 1012.920 1966.720 1019.680 ;
        RECT 1774.720 1011.520 1966.320 1012.920 ;
        RECT 1774.720 1003.400 1966.720 1011.520 ;
        RECT 1775.120 1002.000 1966.720 1003.400 ;
        RECT 1774.720 995.240 1966.720 1002.000 ;
        RECT 1774.720 993.840 1966.320 995.240 ;
      LAYER met3 ;
        RECT 1966.720 994.240 1970.720 994.840 ;
      LAYER met3 ;
        RECT 1774.720 985.720 1966.720 993.840 ;
      LAYER met3 ;
        RECT 1968.190 993.305 1968.490 994.240 ;
        RECT 1968.190 992.990 1968.735 993.305 ;
        RECT 1968.405 992.975 1968.735 992.990 ;
        RECT 1755.630 985.130 1756.010 985.140 ;
        RECT 1770.720 985.130 1774.720 985.320 ;
        RECT 1755.630 984.830 1774.720 985.130 ;
        RECT 1755.630 984.820 1756.010 984.830 ;
        RECT 1770.720 984.720 1774.720 984.830 ;
      LAYER met3 ;
        RECT 1775.120 984.320 1966.720 985.720 ;
        RECT 1774.720 977.560 1966.720 984.320 ;
        RECT 1774.720 976.160 1966.320 977.560 ;
      LAYER met3 ;
        RECT 1966.720 976.560 1970.720 977.160 ;
      LAYER met3 ;
        RECT 1774.720 968.040 1966.720 976.160 ;
      LAYER met3 ;
        RECT 1969.110 974.265 1969.410 976.560 ;
        RECT 1969.110 973.950 1969.655 974.265 ;
        RECT 1969.325 973.935 1969.655 973.950 ;
      LAYER met3 ;
        RECT 1775.120 966.640 1966.720 968.040 ;
        RECT 1774.720 959.880 1966.720 966.640 ;
        RECT 1774.720 958.480 1966.320 959.880 ;
        RECT 1774.720 951.720 1966.720 958.480 ;
        RECT 1775.120 950.320 1966.720 951.720 ;
        RECT 1774.720 943.560 1966.720 950.320 ;
      LAYER met3 ;
        RECT 1968.865 945.010 1969.195 945.025 ;
        RECT 1968.865 944.695 1969.410 945.010 ;
      LAYER met3 ;
        RECT 1774.720 942.160 1966.320 943.560 ;
      LAYER met3 ;
        RECT 1969.110 943.160 1969.410 944.695 ;
        RECT 1966.720 942.560 1970.720 943.160 ;
      LAYER met3 ;
        RECT 1774.720 934.040 1966.720 942.160 ;
      LAYER met3 ;
        RECT 1752.665 933.450 1752.995 933.465 ;
        RECT 1770.720 933.450 1774.720 933.640 ;
        RECT 1752.665 933.150 1774.720 933.450 ;
        RECT 1752.665 933.135 1752.995 933.150 ;
        RECT 1770.720 933.040 1774.720 933.150 ;
      LAYER met3 ;
        RECT 1775.120 932.640 1966.720 934.040 ;
        RECT 1774.720 925.880 1966.720 932.640 ;
        RECT 1774.720 925.015 1966.320 925.880 ;
        RECT 276.000 921.760 1467.600 923.160 ;
      LAYER met3 ;
        RECT 1468.000 922.570 1472.000 922.760 ;
        RECT 1487.245 922.570 1487.575 922.585 ;
        RECT 1468.000 922.270 1487.575 922.570 ;
        RECT 1468.000 922.160 1472.000 922.270 ;
        RECT 1487.245 922.255 1487.575 922.270 ;
      LAYER met3 ;
        RECT 276.000 909.560 1471.730 921.760 ;
      LAYER met3 ;
        RECT 272.000 908.560 276.000 909.160 ;
        RECT 270.750 906.250 271.130 906.260 ;
        RECT 272.630 906.250 272.930 908.560 ;
      LAYER met3 ;
        RECT 276.400 908.160 1471.730 909.560 ;
      LAYER met3 ;
        RECT 270.750 905.950 272.930 906.250 ;
        RECT 270.750 905.940 271.130 905.950 ;
      LAYER met3 ;
        RECT 276.000 745.000 1471.730 908.160 ;
      LAYER met3 ;
        RECT 1484.230 906.250 1484.610 906.260 ;
        RECT 1531.150 906.250 1531.530 906.260 ;
        RECT 1484.230 905.950 1531.530 906.250 ;
        RECT 1484.230 905.940 1484.610 905.950 ;
        RECT 1531.150 905.940 1531.530 905.950 ;
        RECT 1580.830 906.250 1581.210 906.260 ;
        RECT 1627.750 906.250 1628.130 906.260 ;
        RECT 1580.830 905.950 1628.130 906.250 ;
        RECT 1580.830 905.940 1581.210 905.950 ;
        RECT 1627.750 905.940 1628.130 905.950 ;
        RECT 1703.190 906.250 1703.570 906.260 ;
        RECT 1724.350 906.250 1724.730 906.260 ;
        RECT 1703.190 905.950 1724.730 906.250 ;
        RECT 1703.190 905.940 1703.570 905.950 ;
        RECT 1724.350 905.940 1724.730 905.950 ;
        RECT 1773.110 906.250 1773.490 906.260 ;
        RECT 1847.630 906.250 1848.010 906.260 ;
        RECT 1773.110 905.950 1848.010 906.250 ;
        RECT 1773.110 905.940 1773.490 905.950 ;
        RECT 1847.630 905.940 1848.010 905.950 ;
      LAYER met3 ;
        RECT 276.000 743.600 1467.600 745.000 ;
      LAYER met3 ;
        RECT 1468.000 744.410 1472.000 744.600 ;
        RECT 1487.705 744.410 1488.035 744.425 ;
        RECT 1468.000 744.110 1488.035 744.410 ;
        RECT 1468.000 744.000 1472.000 744.110 ;
        RECT 1487.705 744.095 1488.035 744.110 ;
        RECT 272.590 734.580 272.970 734.900 ;
        RECT 272.630 732.360 272.930 734.580 ;
      LAYER met3 ;
        RECT 276.000 732.760 1471.730 743.600 ;
      LAYER met3 ;
        RECT 1579.910 736.250 1580.290 736.260 ;
        RECT 1607.510 736.250 1607.890 736.260 ;
        RECT 1579.910 735.950 1607.890 736.250 ;
        RECT 1579.910 735.940 1580.290 735.950 ;
        RECT 1607.510 735.940 1607.890 735.950 ;
        RECT 272.000 731.760 276.000 732.360 ;
      LAYER met3 ;
        RECT 276.400 731.360 1471.730 732.760 ;
        RECT 276.000 568.200 1471.730 731.360 ;
        RECT 276.000 566.800 1467.600 568.200 ;
      LAYER met3 ;
        RECT 1468.000 567.610 1472.000 567.800 ;
        RECT 1487.245 567.610 1487.575 567.625 ;
        RECT 1468.000 567.310 1487.575 567.610 ;
        RECT 1468.000 567.200 1472.000 567.310 ;
        RECT 1487.245 567.295 1487.575 567.310 ;
      LAYER met3 ;
        RECT 276.000 554.600 1471.730 566.800 ;
      LAYER met3 ;
        RECT 261.805 554.010 262.135 554.025 ;
        RECT 272.000 554.010 276.000 554.200 ;
        RECT 261.805 553.710 276.000 554.010 ;
        RECT 261.805 553.695 262.135 553.710 ;
        RECT 272.000 553.600 276.000 553.710 ;
      LAYER met3 ;
        RECT 276.400 553.200 1471.730 554.600 ;
        RECT 276.000 472.475 1471.730 553.200 ;
      LAYER met3 ;
        RECT 261.805 471.730 262.135 471.745 ;
        RECT 1904.670 471.730 1905.050 471.740 ;
        RECT 261.805 471.430 1905.050 471.730 ;
        RECT 261.805 471.415 262.135 471.430 ;
        RECT 1904.670 471.420 1905.050 471.430 ;
      LAYER via3 ;
        RECT 261.580 1264.980 261.900 1265.300 ;
        RECT 1545.900 1140.540 1546.220 1140.860 ;
        RECT 1592.820 1140.540 1593.140 1140.860 ;
        RECT 1646.180 1140.540 1646.500 1140.860 ;
        RECT 1689.420 1140.540 1689.740 1140.860 ;
        RECT 1739.100 1140.540 1739.420 1140.860 ;
        RECT 1786.020 1140.540 1786.340 1140.860 ;
        RECT 1800.740 1133.740 1801.060 1134.060 ;
        RECT 1783.260 1131.700 1783.580 1132.020 ;
        RECT 1904.700 1118.100 1905.020 1118.420 ;
        RECT 1918.500 1118.100 1918.820 1118.420 ;
        RECT 272.620 1084.100 272.940 1084.420 ;
        RECT 1755.660 984.820 1755.980 985.140 ;
        RECT 270.780 905.940 271.100 906.260 ;
        RECT 1484.260 905.940 1484.580 906.260 ;
        RECT 1531.180 905.940 1531.500 906.260 ;
        RECT 1580.860 905.940 1581.180 906.260 ;
        RECT 1627.780 905.940 1628.100 906.260 ;
        RECT 1703.220 905.940 1703.540 906.260 ;
        RECT 1724.380 905.940 1724.700 906.260 ;
        RECT 1773.140 905.940 1773.460 906.260 ;
        RECT 1847.660 905.940 1847.980 906.260 ;
        RECT 272.620 734.580 272.940 734.900 ;
        RECT 1579.940 735.940 1580.260 736.260 ;
        RECT 1607.540 735.940 1607.860 736.260 ;
        RECT 1904.700 471.420 1905.020 471.740 ;
      LAYER met4 ;
        RECT 261.575 1264.975 261.905 1265.305 ;
        RECT 261.590 1134.490 261.890 1264.975 ;
        RECT 261.150 1133.310 262.330 1134.490 ;
        RECT 272.615 1084.095 272.945 1084.425 ;
        RECT 272.630 1080.090 272.930 1084.095 ;
        RECT 272.190 1078.910 273.370 1080.090 ;
        RECT 270.350 905.510 271.530 906.690 ;
        RECT 277.710 906.250 278.890 906.690 ;
        RECT 289.670 906.250 290.850 906.690 ;
        RECT 277.710 905.950 290.850 906.250 ;
        RECT 277.710 905.510 278.890 905.950 ;
        RECT 289.670 905.510 290.850 905.950 ;
        RECT 272.190 742.310 273.370 743.490 ;
        RECT 272.630 734.905 272.930 742.310 ;
        RECT 272.615 734.575 272.945 734.905 ;
      LAYER met4 ;
        RECT 296.535 472.400 310.020 1449.360 ;
        RECT 313.020 472.400 328.020 1449.360 ;
        RECT 331.020 472.400 364.020 1449.360 ;
        RECT 367.020 472.400 382.020 1449.360 ;
        RECT 385.020 472.400 400.020 1449.360 ;
        RECT 403.020 472.400 418.020 1449.360 ;
        RECT 421.020 472.400 454.020 1449.360 ;
        RECT 457.020 472.400 472.020 1449.360 ;
        RECT 475.020 472.400 490.020 1449.360 ;
        RECT 493.020 472.400 508.020 1449.360 ;
        RECT 511.020 472.400 544.020 1449.360 ;
        RECT 547.020 472.400 562.020 1449.360 ;
        RECT 565.020 472.400 580.020 1449.360 ;
        RECT 583.020 472.400 598.020 1449.360 ;
        RECT 601.020 472.400 634.020 1449.360 ;
        RECT 637.020 472.400 652.020 1449.360 ;
        RECT 655.020 472.400 670.020 1449.360 ;
        RECT 673.020 472.400 688.020 1449.360 ;
        RECT 691.020 472.400 724.020 1449.360 ;
        RECT 727.020 472.400 742.020 1449.360 ;
        RECT 745.020 472.400 760.020 1449.360 ;
        RECT 763.020 472.400 778.020 1449.360 ;
        RECT 781.020 472.400 814.020 1449.360 ;
        RECT 817.020 472.400 832.020 1449.360 ;
        RECT 835.020 472.400 850.020 1449.360 ;
        RECT 853.020 472.400 868.020 1449.360 ;
        RECT 871.020 472.400 904.020 1449.360 ;
        RECT 907.020 472.400 922.020 1449.360 ;
        RECT 925.020 472.400 940.020 1449.360 ;
        RECT 943.020 472.400 958.020 1449.360 ;
        RECT 961.020 472.400 994.020 1449.360 ;
        RECT 997.020 472.400 1012.020 1449.360 ;
        RECT 1015.020 472.400 1030.020 1449.360 ;
        RECT 1033.020 472.400 1048.020 1449.360 ;
        RECT 1051.020 472.400 1084.020 1449.360 ;
        RECT 1087.020 472.400 1102.020 1449.360 ;
        RECT 1105.020 472.400 1120.020 1449.360 ;
        RECT 1123.020 472.400 1138.020 1449.360 ;
        RECT 1141.020 472.400 1174.020 1449.360 ;
        RECT 1177.020 472.400 1192.020 1449.360 ;
        RECT 1195.020 472.400 1210.020 1449.360 ;
        RECT 1213.020 472.400 1228.020 1449.360 ;
        RECT 1231.020 472.400 1264.020 1449.360 ;
        RECT 1267.020 472.400 1282.020 1449.360 ;
        RECT 1285.020 472.400 1300.020 1449.360 ;
        RECT 1303.020 472.400 1318.020 1449.360 ;
        RECT 1321.020 472.400 1354.020 1449.360 ;
        RECT 1357.020 472.400 1372.020 1449.360 ;
        RECT 1375.020 472.400 1390.020 1449.360 ;
        RECT 1393.020 472.400 1408.020 1449.360 ;
        RECT 1411.020 472.400 1444.020 1449.360 ;
        RECT 1447.020 472.400 1448.960 1449.360 ;
      LAYER met4 ;
        RECT 1449.360 472.400 1450.960 1449.360 ;
      LAYER met4 ;
        RECT 1451.360 472.400 1462.020 1449.360 ;
        RECT 1465.020 472.400 1471.705 1449.360 ;
      LAYER met4 ;
        RECT 1545.470 1140.110 1546.650 1141.290 ;
        RECT 1592.815 1140.535 1593.145 1140.865 ;
        RECT 1592.830 1134.490 1593.130 1140.535 ;
        RECT 1645.750 1140.110 1646.930 1141.290 ;
        RECT 1689.415 1140.535 1689.745 1140.865 ;
        RECT 1689.430 1134.490 1689.730 1140.535 ;
        RECT 1738.670 1140.110 1739.850 1141.290 ;
        RECT 1785.590 1140.110 1786.770 1141.290 ;
        RECT 1592.390 1133.310 1593.570 1134.490 ;
        RECT 1688.990 1133.310 1690.170 1134.490 ;
        RECT 1800.310 1133.310 1801.490 1134.490 ;
        RECT 1783.255 1131.695 1783.585 1132.025 ;
        RECT 1773.630 1086.450 1774.810 1086.890 ;
        RECT 1783.270 1086.450 1783.570 1131.695 ;
        RECT 1904.695 1118.095 1905.025 1118.425 ;
        RECT 1918.495 1118.095 1918.825 1118.425 ;
        RECT 1773.630 1086.150 1783.570 1086.450 ;
        RECT 1773.630 1085.710 1774.810 1086.150 ;
        RECT 1755.655 984.815 1755.985 985.145 ;
        RECT 1483.830 905.510 1485.010 906.690 ;
        RECT 1530.750 905.510 1531.930 906.690 ;
        RECT 1580.430 905.510 1581.610 906.690 ;
        RECT 1627.350 905.510 1628.530 906.690 ;
        RECT 1702.790 905.510 1703.970 906.690 ;
        RECT 1723.950 905.510 1725.130 906.690 ;
        RECT 1755.670 736.690 1755.970 984.815 ;
      LAYER met4 ;
        RECT 1794.480 932.080 1804.020 1109.360 ;
        RECT 1807.020 932.080 1822.020 1109.360 ;
        RECT 1825.020 932.080 1840.020 1109.360 ;
        RECT 1843.020 932.080 1858.020 1109.360 ;
        RECT 1861.020 932.080 1870.880 1109.360 ;
      LAYER met4 ;
        RECT 1871.280 932.080 1872.880 1109.360 ;
      LAYER met4 ;
        RECT 1873.280 932.080 1877.505 1109.360 ;
      LAYER met4 ;
        RECT 1772.710 905.510 1773.890 906.690 ;
        RECT 1847.230 905.510 1848.410 906.690 ;
        RECT 1579.510 735.510 1580.690 736.690 ;
        RECT 1607.110 735.510 1608.290 736.690 ;
        RECT 1755.230 735.510 1756.410 736.690 ;
        RECT 1904.710 471.745 1905.010 1118.095 ;
        RECT 1918.510 906.690 1918.810 1118.095 ;
        RECT 1918.070 905.510 1919.250 906.690 ;
        RECT 1904.695 471.415 1905.025 471.745 ;
      LAYER met5 ;
        RECT 301.420 1139.900 1367.460 1141.500 ;
        RECT 301.420 1134.700 303.020 1139.900 ;
        RECT 260.940 1133.100 303.020 1134.700 ;
        RECT 1365.860 1134.700 1367.460 1139.900 ;
        RECT 1412.780 1139.900 1450.260 1141.500 ;
        RECT 1412.780 1134.700 1414.380 1139.900 ;
        RECT 1448.660 1138.100 1450.260 1139.900 ;
        RECT 1509.380 1139.900 1546.860 1141.500 ;
        RECT 1605.980 1139.900 1647.140 1141.500 ;
        RECT 1702.580 1139.900 1740.060 1141.500 ;
        RECT 1785.380 1139.900 1800.780 1141.500 ;
        RECT 1448.660 1136.500 1497.180 1138.100 ;
        RECT 1365.860 1133.100 1414.380 1134.700 ;
        RECT 1495.580 1134.700 1497.180 1136.500 ;
        RECT 1509.380 1134.700 1510.980 1139.900 ;
        RECT 1605.980 1134.700 1607.580 1139.900 ;
        RECT 1702.580 1134.700 1704.180 1139.900 ;
        RECT 1495.580 1133.100 1510.980 1134.700 ;
        RECT 1592.180 1133.100 1607.580 1134.700 ;
        RECT 1688.780 1133.100 1704.180 1134.700 ;
        RECT 1799.180 1134.700 1800.780 1139.900 ;
        RECT 1799.180 1133.100 1801.700 1134.700 ;
        RECT 322.580 1083.700 325.100 1087.100 ;
        RECT 419.180 1083.700 421.700 1087.100 ;
        RECT 515.780 1083.700 518.300 1087.100 ;
        RECT 612.380 1083.700 614.900 1087.100 ;
        RECT 708.980 1083.700 711.500 1087.100 ;
        RECT 805.580 1083.700 808.100 1087.100 ;
        RECT 902.180 1083.700 904.700 1087.100 ;
        RECT 998.780 1083.700 1001.300 1087.100 ;
        RECT 1095.380 1083.700 1097.900 1087.100 ;
        RECT 1191.980 1083.700 1194.500 1087.100 ;
        RECT 1288.580 1083.700 1291.100 1087.100 ;
        RECT 1385.180 1083.700 1387.700 1087.100 ;
        RECT 322.580 1082.100 354.540 1083.700 ;
        RECT 322.580 1080.300 324.180 1082.100 ;
        RECT 271.980 1078.700 324.180 1080.300 ;
        RECT 352.940 1080.300 354.540 1082.100 ;
        RECT 419.180 1082.100 451.140 1083.700 ;
        RECT 419.180 1080.300 420.780 1082.100 ;
        RECT 352.940 1078.700 420.780 1080.300 ;
        RECT 449.540 1080.300 451.140 1082.100 ;
        RECT 515.780 1082.100 547.740 1083.700 ;
        RECT 515.780 1080.300 517.380 1082.100 ;
        RECT 449.540 1078.700 517.380 1080.300 ;
        RECT 546.140 1080.300 547.740 1082.100 ;
        RECT 612.380 1082.100 644.340 1083.700 ;
        RECT 612.380 1080.300 613.980 1082.100 ;
        RECT 546.140 1078.700 613.980 1080.300 ;
        RECT 642.740 1080.300 644.340 1082.100 ;
        RECT 708.980 1082.100 740.940 1083.700 ;
        RECT 708.980 1080.300 710.580 1082.100 ;
        RECT 642.740 1078.700 710.580 1080.300 ;
        RECT 739.340 1080.300 740.940 1082.100 ;
        RECT 805.580 1082.100 837.540 1083.700 ;
        RECT 805.580 1080.300 807.180 1082.100 ;
        RECT 739.340 1078.700 807.180 1080.300 ;
        RECT 835.940 1080.300 837.540 1082.100 ;
        RECT 902.180 1082.100 934.140 1083.700 ;
        RECT 902.180 1080.300 903.780 1082.100 ;
        RECT 835.940 1078.700 903.780 1080.300 ;
        RECT 932.540 1080.300 934.140 1082.100 ;
        RECT 998.780 1082.100 1030.740 1083.700 ;
        RECT 998.780 1080.300 1000.380 1082.100 ;
        RECT 932.540 1078.700 1000.380 1080.300 ;
        RECT 1029.140 1080.300 1030.740 1082.100 ;
        RECT 1095.380 1082.100 1127.340 1083.700 ;
        RECT 1095.380 1080.300 1096.980 1082.100 ;
        RECT 1029.140 1078.700 1096.980 1080.300 ;
        RECT 1125.740 1080.300 1127.340 1082.100 ;
        RECT 1191.980 1082.100 1223.940 1083.700 ;
        RECT 1191.980 1080.300 1193.580 1082.100 ;
        RECT 1125.740 1078.700 1193.580 1080.300 ;
        RECT 1222.340 1080.300 1223.940 1082.100 ;
        RECT 1288.580 1082.100 1320.540 1083.700 ;
        RECT 1288.580 1080.300 1290.180 1082.100 ;
        RECT 1222.340 1078.700 1290.180 1080.300 ;
        RECT 1318.940 1080.300 1320.540 1082.100 ;
        RECT 1385.180 1082.100 1416.220 1083.700 ;
        RECT 1385.180 1080.300 1386.780 1082.100 ;
        RECT 1318.940 1078.700 1386.780 1080.300 ;
        RECT 1414.620 1080.300 1416.220 1082.100 ;
        RECT 1481.780 1080.300 1484.300 1087.100 ;
        RECT 1558.140 1085.500 1580.900 1087.100 ;
        RECT 1558.140 1083.700 1559.740 1085.500 ;
        RECT 1510.300 1082.100 1559.740 1083.700 ;
        RECT 1510.300 1080.300 1511.900 1082.100 ;
        RECT 1414.620 1078.700 1511.900 1080.300 ;
        RECT 1579.300 1080.300 1580.900 1085.500 ;
        RECT 1654.740 1085.500 1677.500 1087.100 ;
        RECT 1654.740 1083.700 1656.340 1085.500 ;
        RECT 1606.900 1082.100 1656.340 1083.700 ;
        RECT 1606.900 1080.300 1608.500 1082.100 ;
        RECT 1579.300 1078.700 1608.500 1080.300 ;
        RECT 1675.900 1080.300 1677.500 1085.500 ;
        RECT 1751.340 1085.500 1775.020 1087.100 ;
        RECT 1751.340 1083.700 1752.940 1085.500 ;
        RECT 1703.500 1082.100 1752.940 1083.700 ;
        RECT 1703.500 1080.300 1705.100 1082.100 ;
        RECT 1675.900 1078.700 1705.100 1080.300 ;
      LAYER met5 ;
        RECT 1132.180 920.300 1145.740 921.900 ;
      LAYER met5 ;
        RECT -768.195 905.300 1485.220 906.900 ;
        RECT 1530.540 905.300 1581.820 906.900 ;
        RECT 1627.140 905.300 1704.180 906.900 ;
        RECT 1723.740 905.300 1774.100 906.900 ;
        RECT 1847.020 905.300 1919.460 906.900 ;
        RECT 271.980 742.100 324.180 743.700 ;
        RECT 322.580 740.300 324.180 742.100 ;
        RECT 352.020 742.100 420.780 743.700 ;
        RECT 352.020 740.300 353.620 742.100 ;
        RECT 322.580 738.700 353.620 740.300 ;
        RECT 419.180 740.300 420.780 742.100 ;
        RECT 448.620 742.100 517.380 743.700 ;
        RECT 448.620 740.300 450.220 742.100 ;
        RECT 419.180 738.700 450.220 740.300 ;
        RECT 515.780 740.300 517.380 742.100 ;
        RECT 545.220 742.100 613.980 743.700 ;
        RECT 545.220 740.300 546.820 742.100 ;
        RECT 515.780 738.700 546.820 740.300 ;
        RECT 612.380 740.300 613.980 742.100 ;
        RECT 641.820 742.100 710.580 743.700 ;
        RECT 641.820 740.300 643.420 742.100 ;
        RECT 612.380 738.700 643.420 740.300 ;
        RECT 708.980 740.300 710.580 742.100 ;
        RECT 738.420 742.100 807.180 743.700 ;
        RECT 738.420 740.300 740.020 742.100 ;
        RECT 708.980 738.700 740.020 740.300 ;
        RECT 805.580 740.300 807.180 742.100 ;
        RECT 835.020 742.100 903.780 743.700 ;
        RECT 835.020 740.300 836.620 742.100 ;
        RECT 805.580 738.700 836.620 740.300 ;
        RECT 902.180 740.300 903.780 742.100 ;
        RECT 931.620 742.100 1000.380 743.700 ;
        RECT 931.620 740.300 933.220 742.100 ;
        RECT 902.180 738.700 933.220 740.300 ;
        RECT 998.780 740.300 1000.380 742.100 ;
        RECT 1028.220 742.100 1096.980 743.700 ;
        RECT 1028.220 740.300 1029.820 742.100 ;
        RECT 998.780 738.700 1029.820 740.300 ;
        RECT 1095.380 740.300 1096.980 742.100 ;
        RECT 1124.820 742.100 1193.580 743.700 ;
        RECT 1124.820 740.300 1126.420 742.100 ;
        RECT 1095.380 738.700 1126.420 740.300 ;
        RECT 1191.980 740.300 1193.580 742.100 ;
        RECT 1221.420 742.100 1290.180 743.700 ;
        RECT 1221.420 740.300 1223.020 742.100 ;
        RECT 1191.980 738.700 1223.020 740.300 ;
        RECT 1288.580 740.300 1290.180 742.100 ;
        RECT 1318.020 742.100 1386.780 743.700 ;
        RECT 1318.020 740.300 1319.620 742.100 ;
        RECT 1288.580 738.700 1319.620 740.300 ;
        RECT 1385.180 740.300 1386.780 742.100 ;
        RECT 1414.620 742.100 1478.780 743.700 ;
        RECT 1414.620 740.300 1416.220 742.100 ;
        RECT 1385.180 738.700 1416.220 740.300 ;
        RECT 322.580 735.300 325.100 738.700 ;
        RECT 419.180 735.300 421.700 738.700 ;
        RECT 515.780 735.300 518.300 738.700 ;
        RECT 612.380 735.300 614.900 738.700 ;
        RECT 708.980 735.300 711.500 738.700 ;
        RECT 805.580 735.300 808.100 738.700 ;
        RECT 902.180 735.300 904.700 738.700 ;
        RECT 998.780 735.300 1001.300 738.700 ;
        RECT 1095.380 735.300 1097.900 738.700 ;
        RECT 1191.980 735.300 1194.500 738.700 ;
        RECT 1288.580 735.300 1291.100 738.700 ;
        RECT 1385.180 735.300 1387.700 738.700 ;
        RECT 1477.180 736.900 1478.780 742.100 ;
        RECT 1488.220 742.100 1532.140 743.700 ;
        RECT 1488.220 736.900 1489.820 742.100 ;
        RECT 1477.180 735.300 1489.820 736.900 ;
        RECT 1530.540 736.900 1532.140 742.100 ;
        RECT 1675.900 742.100 1725.340 743.700 ;
        RECT 1675.900 736.900 1677.500 742.100 ;
        RECT 1530.540 735.300 1580.900 736.900 ;
        RECT 1606.900 735.300 1677.500 736.900 ;
        RECT 1723.740 736.900 1725.340 742.100 ;
        RECT 1723.740 735.300 1756.620 736.900 ;
  END
END user_project_wrapper
END LIBRARY

