VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO decred_hash_macro
  CLASS BLOCK ;
  FOREIGN decred_hash_macro ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 1000.000 ;
  PIN CLK
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 655.130 996.000 655.410 1000.000 ;
    END
  END CLK
  PIN DATA_AVAILABLE
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 724.130 0.000 724.410 4.000 ;
    END
  END DATA_AVAILABLE
  PIN DATA_FROM_HASH[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END DATA_FROM_HASH[0]
  PIN DATA_FROM_HASH[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END DATA_FROM_HASH[1]
  PIN DATA_FROM_HASH[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 896.170 996.000 896.450 1000.000 ;
    END
  END DATA_FROM_HASH[2]
  PIN DATA_FROM_HASH[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1084.770 0.000 1085.050 4.000 ;
    END
  END DATA_FROM_HASH[3]
  PIN DATA_FROM_HASH[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 194.520 1200.000 195.120 ;
    END
  END DATA_FROM_HASH[4]
  PIN DATA_FROM_HASH[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END DATA_FROM_HASH[5]
  PIN DATA_FROM_HASH[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 173.970 996.000 174.250 1000.000 ;
    END
  END DATA_FROM_HASH[6]
  PIN DATA_FROM_HASH[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 715.400 4.000 716.000 ;
    END
  END DATA_FROM_HASH[7]
  PIN DATA_TO_HASH[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 414.090 996.000 414.370 1000.000 ;
    END
  END DATA_TO_HASH[0]
  PIN DATA_TO_HASH[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END DATA_TO_HASH[1]
  PIN DATA_TO_HASH[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 372.680 1200.000 373.280 ;
    END
  END DATA_TO_HASH[2]
  PIN DATA_TO_HASH[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 16.360 1200.000 16.960 ;
    END
  END DATA_TO_HASH[3]
  PIN DATA_TO_HASH[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.200 4.000 892.800 ;
    END
  END DATA_TO_HASH[4]
  PIN DATA_TO_HASH[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END DATA_TO_HASH[5]
  PIN DATA_TO_HASH[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1015.770 996.000 1016.050 1000.000 ;
    END
  END DATA_TO_HASH[6]
  PIN DATA_TO_HASH[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 294.490 996.000 294.770 1000.000 ;
    END
  END DATA_TO_HASH[7]
  PIN HASH_ADDR[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.650 996.000 775.930 1000.000 ;
    END
  END HASH_ADDR[0]
  PIN HASH_ADDR[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.450 996.000 53.730 1000.000 ;
    END
  END HASH_ADDR[1]
  PIN HASH_ADDR[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1136.290 996.000 1136.570 1000.000 ;
    END
  END HASH_ADDR[2]
  PIN HASH_ADDR[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.170 0.000 965.450 4.000 ;
    END
  END HASH_ADDR[3]
  PIN HASH_ADDR[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END HASH_ADDR[4]
  PIN HASH_ADDR[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 905.800 1200.000 906.400 ;
    END
  END HASH_ADDR[5]
  PIN HASH_EN
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 4.000 ;
    END
  END HASH_EN
  PIN MACRO_RD_SELECT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 603.610 0.000 603.890 4.000 ;
    END
  END MACRO_RD_SELECT
  PIN MACRO_WR_SELECT
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 550.840 1200.000 551.440 ;
    END
  END MACRO_WR_SELECT
  PIN THREAD_COUNT[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 727.640 1200.000 728.240 ;
    END
  END THREAD_COUNT[0]
  PIN THREAD_COUNT[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END THREAD_COUNT[1]
  PIN THREAD_COUNT[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 534.610 996.000 534.890 1000.000 ;
    END
  END THREAD_COUNT[2]
  PIN THREAD_COUNT[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 844.650 0.000 844.930 4.000 ;
    END
  END THREAD_COUNT[3]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 987.600 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 987.600 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1194.160 987.445 ;
      LAYER met1 ;
        RECT 3.750 8.540 1194.160 987.600 ;
      LAYER met2 ;
        RECT 1.930 995.720 53.170 996.000 ;
        RECT 54.010 995.720 173.690 996.000 ;
        RECT 174.530 995.720 294.210 996.000 ;
        RECT 295.050 995.720 413.810 996.000 ;
        RECT 414.650 995.720 534.330 996.000 ;
        RECT 535.170 995.720 654.850 996.000 ;
        RECT 655.690 995.720 775.370 996.000 ;
        RECT 776.210 995.720 895.890 996.000 ;
        RECT 896.730 995.720 1015.490 996.000 ;
        RECT 1016.330 995.720 1136.010 996.000 ;
        RECT 1136.850 995.720 1191.300 996.000 ;
        RECT 1.930 4.280 1191.300 995.720 ;
        RECT 1.930 4.000 2.570 4.280 ;
        RECT 3.410 4.000 122.170 4.280 ;
        RECT 123.010 4.000 242.690 4.280 ;
        RECT 243.530 4.000 363.210 4.280 ;
        RECT 364.050 4.000 483.730 4.280 ;
        RECT 484.570 4.000 603.330 4.280 ;
        RECT 604.170 4.000 723.850 4.280 ;
        RECT 724.690 4.000 844.370 4.280 ;
        RECT 845.210 4.000 964.890 4.280 ;
        RECT 965.730 4.000 1084.490 4.280 ;
        RECT 1085.330 4.000 1191.300 4.280 ;
      LAYER met3 ;
        RECT 0.270 906.800 1196.000 987.525 ;
        RECT 0.270 905.400 1195.600 906.800 ;
        RECT 0.270 893.200 1196.000 905.400 ;
        RECT 4.400 891.800 1196.000 893.200 ;
        RECT 0.270 728.640 1196.000 891.800 ;
        RECT 0.270 727.240 1195.600 728.640 ;
        RECT 0.270 716.400 1196.000 727.240 ;
        RECT 4.400 715.000 1196.000 716.400 ;
        RECT 0.270 551.840 1196.000 715.000 ;
        RECT 0.270 550.440 1195.600 551.840 ;
        RECT 0.270 538.240 1196.000 550.440 ;
        RECT 4.400 536.840 1196.000 538.240 ;
        RECT 0.270 373.680 1196.000 536.840 ;
        RECT 0.270 372.280 1195.600 373.680 ;
        RECT 0.270 360.080 1196.000 372.280 ;
        RECT 4.400 358.680 1196.000 360.080 ;
        RECT 0.270 195.520 1196.000 358.680 ;
        RECT 0.270 194.120 1195.600 195.520 ;
        RECT 0.270 181.920 1196.000 194.120 ;
        RECT 4.400 180.520 1196.000 181.920 ;
        RECT 0.270 17.360 1196.000 180.520 ;
        RECT 0.270 15.960 1195.600 17.360 ;
        RECT 0.270 10.715 1196.000 15.960 ;
      LAYER met4 ;
        RECT 0.295 10.640 20.640 987.600 ;
        RECT 23.040 10.640 97.440 987.600 ;
        RECT 99.840 10.640 1175.465 987.600 ;
      LAYER met5 ;
        RECT 326.260 538.100 339.820 539.700 ;
  END
END decred_hash_macro
END LIBRARY

