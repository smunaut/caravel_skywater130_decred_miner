* NGSPICE file created from decred_controller.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

.subckt decred_controller CLK_LED DATA_AVAILABLE DATA_FROM_HASH[0] DATA_FROM_HASH[1]
+ DATA_FROM_HASH[2] DATA_FROM_HASH[3] DATA_FROM_HASH[4] DATA_FROM_HASH[5] DATA_FROM_HASH[6]
+ DATA_FROM_HASH[7] DATA_TO_HASH[0] DATA_TO_HASH[1] DATA_TO_HASH[2] DATA_TO_HASH[3]
+ DATA_TO_HASH[4] DATA_TO_HASH[5] DATA_TO_HASH[6] DATA_TO_HASH[7] EXT_RESET_N_fromHost
+ EXT_RESET_N_toClient HASH_ADDR[0] HASH_ADDR[1] HASH_ADDR[2] HASH_ADDR[3] HASH_ADDR[4]
+ HASH_ADDR[5] HASH_EN HASH_LED ID_fromClient ID_toHost IRQ_OUT_fromClient IRQ_OUT_toHost
+ M1_CLK_IN M1_CLK_SELECT MACRO_RD_SELECT MACRO_WR_SELECT MISO_fromClient MISO_toHost
+ MOSI_fromHost MOSI_toClient PLL_INPUT S1_CLK_IN S1_CLK_SELECT SCLK_fromHost SCLK_toClient
+ SCSN_fromHost SCSN_toClient SPI_CLK_RESET_N THREAD_COUNT[0] THREAD_COUNT[1] THREAD_COUNT[2]
+ THREAD_COUNT[3] m1_clk_local VPWR VGND
X_2106_ _2121_/CLK _1850_/Y VGND VGND VPWR VPWR _1211_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_39_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2037_ _2022_/CLK _1879_/C VGND VGND VPWR VPWR _2031_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_18_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1270_ _1209_/A VGND VGND VPWR VPWR _1365_/A sky130_fd_sc_hd__inv_2
XFILLER_36_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1606_ _1596_/A _1596_/B _1605_/Y VGND VGND VPWR VPWR _1606_/X sky130_fd_sc_hd__o21a_4
X_1468_ _1464_/X _1467_/X _1175_/X VGND VGND VPWR VPWR _1468_/Y sky130_fd_sc_hd__a21oi_4
X_1399_ THREAD_COUNT[2] _1345_/X _1397_/Y _1398_/Y VGND VGND VPWR VPWR _1399_/Y sky130_fd_sc_hd__a22oi_4
X_1537_ _2196_/Q _1525_/X _1536_/X VGND VGND VPWR VPWR _1537_/X sky130_fd_sc_hd__o21a_4
XFILLER_35_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1253_ _1253_/A _1230_/B VGND VGND VPWR VPWR _1253_/Y sky130_fd_sc_hd__nand2_4
X_1322_ _1321_/X VGND VGND VPWR VPWR _1323_/C sky130_fd_sc_hd__buf_2
Xclkbuf_1_0_0_m1_clk_local clkbuf_0_m1_clk_local/X VGND VGND VPWR VPWR clkbuf_2_1_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1184_ _1184_/A _2220_/Q _1184_/C VGND VGND VPWR VPWR _1185_/A sky130_fd_sc_hd__nor3_4
XFILLER_32_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1940_ _1940_/A VGND VGND VPWR VPWR _1940_/Y sky130_fd_sc_hd__inv_2
X_1871_ _1864_/Y VGND VGND VPWR VPWR _1874_/A sky130_fd_sc_hd__buf_2
XFILLER_9_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1236_ _2089_/Q VGND VGND VPWR VPWR _1236_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_0_m1_clk_local m1_clk_local VGND VGND VPWR VPWR clkbuf_0_m1_clk_local/X sky130_fd_sc_hd__clkbuf_16
X_1305_ _1917_/A VGND VGND VPWR VPWR _1307_/B sky130_fd_sc_hd__buf_2
XFILLER_52_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1167_ _1164_/X _2074_/Q _1166_/X VGND VGND VPWR VPWR _1167_/Y sky130_fd_sc_hd__a21oi_4
X_1098_ _1038_/X VGND VGND VPWR VPWR _1446_/A sky130_fd_sc_hd__buf_2
XFILLER_55_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2070_ _2056_/CLK _2070_/D VGND VGND VPWR VPWR _2070_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_3_3_0_m1_clk_local clkbuf_3_3_0_m1_clk_local/A VGND VGND VPWR VPWR _2016_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1021_ _1024_/A _1034_/A _1020_/X VGND VGND VPWR VPWR _1021_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_19_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1785_ _1814_/A _2121_/Q VGND VGND VPWR VPWR _1785_/Y sky130_fd_sc_hd__nand2_4
X_1923_ _1902_/Y _1918_/A _1922_/Y VGND VGND VPWR VPWR _1923_/Y sky130_fd_sc_hd__o21ai_4
X_1854_ _1856_/A _1856_/B VGND VGND VPWR VPWR _1854_/Y sky130_fd_sc_hd__nor2_4
X_1219_ _1312_/A _1218_/X VGND VGND VPWR VPWR _1708_/C sky130_fd_sc_hd__nor2_4
XFILLER_25_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2199_ _2207_/CLK _1532_/X VGND VGND VPWR VPWR _2199_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1570_ _1570_/A SPI_CLK_RESET_N _1570_/C _1569_/X VGND VGND VPWR VPWR _2187_/D sky130_fd_sc_hd__and4_4
XFILLER_3_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2122_ _2127_/CLK _2122_/D VGND VGND VPWR VPWR _1814_/A sky130_fd_sc_hd__dfxtp_4
X_2053_ _2056_/CLK DATA_FROM_HASH[2] VGND VGND VPWR VPWR _2053_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1004_ _1004_/A VGND VGND VPWR VPWR _1004_/X sky130_fd_sc_hd__buf_2
X_1837_ _2113_/Q _1836_/Y VGND VGND VPWR VPWR _1837_/Y sky130_fd_sc_hd__xnor2_4
X_1906_ _1904_/Y _1473_/B _1905_/X _1407_/Y _1889_/X VGND VGND VPWR VPWR _1906_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1768_ _1746_/A _1940_/A _1767_/Y VGND VGND VPWR VPWR _1768_/Y sky130_fd_sc_hd__o21ai_4
X_1699_ _1697_/A _2147_/Q VGND VGND VPWR VPWR _2148_/D sky130_fd_sc_hd__and2_4
XFILLER_25_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1622_ _1621_/C _1609_/A _1609_/C _1609_/D _1101_/X VGND VGND VPWR VPWR _1622_/Y
+ sky130_fd_sc_hd__a41oi_4
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1484_ _1484_/A _2065_/Q VGND VGND VPWR VPWR _1484_/X sky130_fd_sc_hd__xor2_4
X_1553_ _1456_/B VGND VGND VPWR VPWR _1553_/Y sky130_fd_sc_hd__inv_2
X_2036_ _2022_/CLK _2036_/D VGND VGND VPWR VPWR _2036_/Q sky130_fd_sc_hd__dfxtp_4
X_2105_ _2121_/CLK _2105_/D VGND VGND VPWR VPWR _1829_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1605_ _1574_/A _1604_/Y _1599_/X _1596_/A _1101_/X VGND VGND VPWR VPWR _1605_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1536_ _2197_/Q _1526_/X _1535_/X VGND VGND VPWR VPWR _1536_/X sky130_fd_sc_hd__o21a_4
XFILLER_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1467_ _1999_/D _1355_/X _1172_/X _1466_/Y VGND VGND VPWR VPWR _1467_/X sky130_fd_sc_hd__a211o_4
X_1398_ _2101_/Q _1397_/B _1708_/C _1708_/A VGND VGND VPWR VPWR _1398_/Y sky130_fd_sc_hd__a2bb2oi_4
X_2019_ _2110_/CLK _2019_/D VGND VGND VPWR VPWR DATA_TO_HASH[0] sky130_fd_sc_hd__dfxtp_4
XFILLER_50_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1252_ _1252_/A _1252_/B VGND VGND VPWR VPWR _1252_/Y sky130_fd_sc_hd__nand2_4
X_1321_ _1971_/A _1320_/Y _1066_/A _1066_/D _1001_/A VGND VGND VPWR VPWR _1321_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_64_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1183_ _1205_/A VGND VGND VPWR VPWR _1184_/C sky130_fd_sc_hd__inv_2
Xclkbuf_3_4_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_4_9_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_59_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1519_ _1503_/A _1762_/C _1510_/X VGND VGND VPWR VPWR _1519_/X sky130_fd_sc_hd__o21a_4
XFILLER_55_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1870_ _1930_/A _1865_/X _1869_/Y VGND VGND VPWR VPWR _2097_/D sky130_fd_sc_hd__o21ai_4
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1235_ _1232_/Y _1233_/X _1234_/Y VGND VGND VPWR VPWR _1235_/Y sky130_fd_sc_hd__o21ai_4
X_1166_ _1166_/A VGND VGND VPWR VPWR _1166_/X sky130_fd_sc_hd__buf_2
X_1304_ _1863_/B VGND VGND VPWR VPWR _1917_/A sky130_fd_sc_hd__buf_2
X_1097_ _1058_/A VGND VGND VPWR VPWR _1097_/Y sky130_fd_sc_hd__inv_2
X_1999_ _2127_/CLK _1999_/D VGND VGND VPWR VPWR _1999_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_47_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1020_ _2242_/Q _1016_/B VGND VGND VPWR VPWR _1020_/X sky130_fd_sc_hd__or2_4
X_1922_ _1924_/A _1918_/B _1922_/C VGND VGND VPWR VPWR _1922_/Y sky130_fd_sc_hd__nand3_4
XFILLER_34_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1784_ _1784_/A VGND VGND VPWR VPWR _1813_/D sky130_fd_sc_hd__inv_2
X_1853_ _1772_/A _1852_/Y VGND VGND VPWR VPWR _2104_/D sky130_fd_sc_hd__xor2_4
XFILLER_29_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1218_ _1184_/C VGND VGND VPWR VPWR _1218_/X sky130_fd_sc_hd__buf_2
X_1149_ _1149_/A _1149_/B VGND VGND VPWR VPWR _1150_/A sky130_fd_sc_hd__nor2_4
X_2198_ _2207_/CLK _1534_/X VGND VGND VPWR VPWR _2198_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_52_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2121_ _2121_/CLK _1816_/X VGND VGND VPWR VPWR _2121_/Q sky130_fd_sc_hd__dfxtp_4
X_2052_ _2083_/CLK DATA_FROM_HASH[1] VGND VGND VPWR VPWR _2044_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_19_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1003_ _1003_/A VGND VGND VPWR VPWR _1003_/X sky130_fd_sc_hd__buf_2
X_1905_ _1905_/A VGND VGND VPWR VPWR _1905_/X sky130_fd_sc_hd__buf_2
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1836_ _1836_/A _1836_/B _1836_/C _1831_/Y VGND VGND VPWR VPWR _1836_/Y sky130_fd_sc_hd__nand4_4
X_1767_ _1739_/A _1867_/B _2131_/Q VGND VGND VPWR VPWR _1767_/Y sky130_fd_sc_hd__nand3_4
X_1698_ _1697_/A SCLK_fromHost VGND VGND VPWR VPWR _1698_/X sky130_fd_sc_hd__and2_4
XFILLER_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1621_ _1619_/Y _1621_/B _1621_/C _1609_/D VGND VGND VPWR VPWR _1621_/X sky130_fd_sc_hd__and4_4
X_1552_ _1551_/X VGND VGND VPWR VPWR _1552_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2104_ _2110_/CLK _2104_/D VGND VGND VPWR VPWR _1772_/A sky130_fd_sc_hd__dfxtp_4
X_1483_ _1105_/B _2059_/Q VGND VGND VPWR VPWR _1483_/X sky130_fd_sc_hd__xor2_4
XFILLER_62_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2035_ _2027_/CLK _1883_/C VGND VGND VPWR VPWR _2029_/D sky130_fd_sc_hd__dfxtp_4
X_1819_ _1827_/B _1813_/C VGND VGND VPWR VPWR _1820_/B sky130_fd_sc_hd__nand2_4
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1604_ _1595_/C VGND VGND VPWR VPWR _1604_/Y sky130_fd_sc_hd__inv_2
X_1535_ _1504_/A VGND VGND VPWR VPWR _1535_/X sky130_fd_sc_hd__buf_2
X_1397_ _1395_/Y _1397_/B _1396_/Y VGND VGND VPWR VPWR _1397_/Y sky130_fd_sc_hd__nand3_4
X_1466_ _1387_/X _1466_/B VGND VGND VPWR VPWR _1466_/Y sky130_fd_sc_hd__nor2_4
XFILLER_50_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2018_ _2181_/CLK _2131_/Q VGND VGND VPWR VPWR _2017_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1320_ _1309_/A VGND VGND VPWR VPWR _1320_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1182_ _1148_/A _1150_/A _1048_/A VGND VGND VPWR VPWR _1189_/A sky130_fd_sc_hd__nand3_4
X_1251_ _1274_/A _1251_/B VGND VGND VPWR VPWR _1252_/B sky130_fd_sc_hd__nand2_4
XFILLER_64_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1449_ _1449_/A _1309_/A _1449_/C VGND VGND VPWR VPWR _1449_/Y sky130_fd_sc_hd__nor3_4
X_1518_ _1501_/Y _2196_/Q _1517_/X VGND VGND VPWR VPWR _1518_/X sky130_fd_sc_hd__o21a_4
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1303_ _1753_/C _1279_/Y _1283_/A _1302_/Y VGND VGND VPWR VPWR _1307_/A sky130_fd_sc_hd__a211o_4
XFILLER_49_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1234_ _1164_/X _2073_/Q _1166_/A VGND VGND VPWR VPWR _1234_/Y sky130_fd_sc_hd__a21oi_4
X_1165_ _1172_/A VGND VGND VPWR VPWR _1166_/A sky130_fd_sc_hd__inv_2
XFILLER_37_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1096_ _1894_/A _1966_/B _1079_/X VGND VGND VPWR VPWR _1096_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_20_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1998_ _2022_/CLK _2086_/Q VGND VGND VPWR VPWR _1998_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_28_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1921_ _1316_/Y _1918_/A _1920_/Y VGND VGND VPWR VPWR _1921_/Y sky130_fd_sc_hd__o21ai_4
X_1852_ _1477_/Y _1856_/A _1856_/B VGND VGND VPWR VPWR _1852_/Y sky130_fd_sc_hd__nor3_4
X_1783_ _1783_/A _1817_/B VGND VGND VPWR VPWR _1784_/A sky130_fd_sc_hd__nand2_4
XFILLER_6_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1217_ _1145_/A VGND VGND VPWR VPWR _1217_/X sky130_fd_sc_hd__buf_2
X_1148_ _1148_/A VGND VGND VPWR VPWR _1207_/C sky130_fd_sc_hd__buf_2
X_2197_ _2207_/CLK _1537_/X VGND VGND VPWR VPWR _2197_/Q sky130_fd_sc_hd__dfxtp_4
X_1079_ _1067_/Y VGND VGND VPWR VPWR _1079_/X sky130_fd_sc_hd__buf_2
XFILLER_52_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2120_ _2121_/CLK _1818_/Y VGND VGND VPWR VPWR _1783_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_39_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2051_ _2042_/CLK DATA_FROM_HASH[0] VGND VGND VPWR VPWR _2043_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1002_ _1004_/A VGND VGND VPWR VPWR _1003_/A sky130_fd_sc_hd__buf_2
X_1835_ _1834_/X VGND VGND VPWR VPWR _1836_/A sky130_fd_sc_hd__buf_2
X_1904_ _1904_/A VGND VGND VPWR VPWR _1904_/Y sky130_fd_sc_hd__inv_2
X_1766_ _1750_/A VGND VGND VPWR VPWR _1867_/B sky130_fd_sc_hd__buf_2
X_1697_ _1697_/A _2149_/Q VGND VGND VPWR VPWR _2150_/D sky130_fd_sc_hd__and2_4
XFILLER_40_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1482_ _2060_/Q _1482_/B VGND VGND VPWR VPWR _1482_/Y sky130_fd_sc_hd__nor2_4
X_1620_ _1576_/A VGND VGND VPWR VPWR _1621_/B sky130_fd_sc_hd__buf_2
X_1551_ _1545_/B _1549_/Y _1550_/Y VGND VGND VPWR VPWR _1551_/X sky130_fd_sc_hd__a21o_4
XFILLER_8_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2103_ _2110_/CLK _1855_/X VGND VGND VPWR VPWR _2103_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2034_ _2181_/CLK _2034_/D VGND VGND VPWR VPWR HASH_ADDR[5] sky130_fd_sc_hd__dfxtp_4
X_1818_ _1783_/A _1818_/B VGND VGND VPWR VPWR _1818_/Y sky130_fd_sc_hd__xnor2_4
X_1749_ _1739_/A VGND VGND VPWR VPWR _1763_/A sky130_fd_sc_hd__buf_2
XFILLER_45_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_4_0_addressalyzerBlock.SPI_CLK clkbuf_3_2_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2083_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_42_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1465_ _2039_/D VGND VGND VPWR VPWR _1466_/B sky130_fd_sc_hd__inv_2
X_1603_ _1596_/C _1601_/Y _1602_/Y VGND VGND VPWR VPWR _1603_/X sky130_fd_sc_hd__o21a_4
X_1534_ _2197_/Q _1525_/X _1533_/X VGND VGND VPWR VPWR _1534_/X sky130_fd_sc_hd__o21a_4
X_1396_ _1419_/A _2109_/Q _1419_/C VGND VGND VPWR VPWR _1396_/Y sky130_fd_sc_hd__nand3_4
X_2017_ _2181_/CLK _2017_/D VGND VGND VPWR VPWR MACRO_WR_SELECT sky130_fd_sc_hd__dfxtp_4
XFILLER_35_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1181_ _1088_/X _1177_/Y _1180_/X VGND VGND VPWR VPWR _1181_/Y sky130_fd_sc_hd__o21ai_4
X_1250_ _1246_/Y _1247_/Y _1249_/X VGND VGND VPWR VPWR _1252_/A sky130_fd_sc_hd__a21o_4
XFILLER_32_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1517_ _1503_/A _1902_/A _1510_/X VGND VGND VPWR VPWR _1517_/X sky130_fd_sc_hd__o21a_4
X_1448_ _1438_/A _1451_/B _1451_/C VGND VGND VPWR VPWR _1448_/Y sky130_fd_sc_hd__nor3_4
XFILLER_55_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1379_ _2077_/Q VGND VGND VPWR VPWR _1922_/C sky130_fd_sc_hd__buf_2
XFILLER_11_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1233_ _1170_/A VGND VGND VPWR VPWR _1233_/X sky130_fd_sc_hd__buf_2
X_1302_ _1086_/X _1049_/X _1296_/Y VGND VGND VPWR VPWR _1302_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_52_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1164_ _1170_/A VGND VGND VPWR VPWR _1164_/X sky130_fd_sc_hd__buf_2
XFILLER_37_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1095_ _1748_/C VGND VGND VPWR VPWR _1894_/A sky130_fd_sc_hd__buf_2
X_1997_ _2027_/CLK _2085_/Q VGND VGND VPWR VPWR _1997_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_20_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0_addressalyzerBlock.SPI_CLK clkbuf_0_addressalyzerBlock.SPI_CLK/X VGND
+ VGND VPWR VPWR clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_7_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1851_ _1829_/C _1851_/B VGND VGND VPWR VPWR _2105_/D sky130_fd_sc_hd__xor2_4
X_1920_ _1924_/A _1918_/B HASH_LED VGND VGND VPWR VPWR _1920_/Y sky130_fd_sc_hd__nand3_4
X_1782_ _1782_/A VGND VGND VPWR VPWR _1813_/C sky130_fd_sc_hd__buf_2
X_1216_ _1216_/A _1215_/Y VGND VGND VPWR VPWR _1223_/A sky130_fd_sc_hd__nor2_4
XFILLER_29_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2196_ _2207_/CLK _1539_/X VGND VGND VPWR VPWR _2196_/Q sky130_fd_sc_hd__dfxtp_4
X_1147_ _1147_/A _1147_/B VGND VGND VPWR VPWR _1148_/A sky130_fd_sc_hd__nor2_4
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1078_ _1278_/B VGND VGND VPWR VPWR _1966_/B sky130_fd_sc_hd__buf_2
XFILLER_29_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2050_ _2050_/CLK _2050_/D VGND VGND VPWR VPWR _1180_/A sky130_fd_sc_hd__dfxtp_4
X_1001_ _1001_/A VGND VGND VPWR VPWR _1004_/A sky130_fd_sc_hd__inv_2
XFILLER_15_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1903_ _1902_/Y _1885_/X _1888_/X _1383_/Y _1890_/X VGND VGND VPWR VPWR _1903_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1834_ _1851_/B _1829_/B _1829_/C VGND VGND VPWR VPWR _1834_/X sky130_fd_sc_hd__and3_4
X_1765_ _1633_/A _1740_/X _1139_/A VGND VGND VPWR VPWR _1940_/A sky130_fd_sc_hd__nand3_4
X_1696_ _1696_/A SCSN_fromHost VGND VGND VPWR VPWR _2151_/D sky130_fd_sc_hd__or2_4
XFILLER_57_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2179_ _2181_/CLK _2179_/D VGND VGND VPWR VPWR _1587_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_15_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1481_ _1479_/X _1223_/A _1480_/X VGND VGND VPWR VPWR _2212_/D sky130_fd_sc_hd__a21o_4
X_1550_ _1545_/B _1549_/Y _1457_/A VGND VGND VPWR VPWR _1550_/Y sky130_fd_sc_hd__o21ai_4
X_2033_ _2127_/CLK _2039_/Q VGND VGND VPWR VPWR HASH_ADDR[4] sky130_fd_sc_hd__dfxtp_4
X_2102_ _2110_/CLK _2102_/D VGND VGND VPWR VPWR _2102_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1817_ _1827_/B _1817_/B _1813_/C VGND VGND VPWR VPWR _1818_/B sky130_fd_sc_hd__nand3_4
X_1748_ _1633_/A _1740_/X _1748_/C VGND VGND VPWR VPWR _1932_/A sky130_fd_sc_hd__nand3_4
X_1679_ _2160_/Q VGND VGND VPWR VPWR _1693_/B sky130_fd_sc_hd__inv_2
XFILLER_42_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1602_ _1599_/X _1600_/A _1596_/A _1596_/C _1101_/X VGND VGND VPWR VPWR _1602_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1395_ _1378_/Y _1393_/Y _1394_/X VGND VGND VPWR VPWR _1395_/Y sky130_fd_sc_hd__o21ai_4
X_1464_ _1918_/C _1355_/X _1166_/X _1463_/Y VGND VGND VPWR VPWR _1464_/X sky130_fd_sc_hd__a211o_4
X_1533_ _2198_/Q _1526_/X _1521_/X VGND VGND VPWR VPWR _1533_/X sky130_fd_sc_hd__o21a_4
X_2016_ _2016_/CLK _2015_/Q VGND VGND VPWR VPWR HASH_EN sky130_fd_sc_hd__dfxtp_4
XFILLER_50_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1180_ _1180_/A _1180_/B VGND VGND VPWR VPWR _1180_/X sky130_fd_sc_hd__or2_4
XFILLER_49_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1516_ _1501_/Y _2197_/Q _1515_/X VGND VGND VPWR VPWR _2205_/D sky130_fd_sc_hd__o21a_4
XFILLER_59_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1378_ _1788_/A _1265_/B _1732_/A _1473_/B _1473_/C VGND VGND VPWR VPWR _1378_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1447_ _1441_/Y _1445_/Y _1446_/X VGND VGND VPWR VPWR _1447_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1232_ _1232_/A VGND VGND VPWR VPWR _1232_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1301_ _1297_/X _1300_/X _1040_/X VGND VGND VPWR VPWR _2225_/D sky130_fd_sc_hd__a21oi_4
XFILLER_64_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1163_ _2082_/Q VGND VGND VPWR VPWR _1163_/Y sky130_fd_sc_hd__inv_2
X_1094_ _1058_/X _1090_/X _1093_/Y VGND VGND VPWR VPWR _1094_/Y sky130_fd_sc_hd__o21ai_4
X_1996_ _2016_/CLK _2084_/Q VGND VGND VPWR VPWR _1996_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1781_ _1781_/A _2117_/Q _2116_/Q _2115_/Q VGND VGND VPWR VPWR _1782_/A sky130_fd_sc_hd__and4_4
X_1850_ _1850_/A VGND VGND VPWR VPWR _1850_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1215_ _1215_/A _1215_/B _1191_/A VGND VGND VPWR VPWR _1215_/Y sky130_fd_sc_hd__nor3_4
X_1146_ _1048_/A VGND VGND VPWR VPWR _1215_/A sky130_fd_sc_hd__buf_2
XFILLER_1_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2195_ _2202_/CLK _1541_/X VGND VGND VPWR VPWR _2195_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1077_ _1484_/A _1076_/X _1072_/Y VGND VGND VPWR VPWR _1077_/Y sky130_fd_sc_hd__o21ai_4
X_1979_ PLL_INPUT M1_CLK_SELECT _1978_/Y VGND VGND VPWR VPWR m1_clk_local sky130_fd_sc_hd__o21a_4
XFILLER_20_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1000_ _1280_/A VGND VGND VPWR VPWR _1001_/A sky130_fd_sc_hd__buf_2
X_1902_ _1902_/A VGND VGND VPWR VPWR _1902_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1833_ _1833_/A _1832_/Y VGND VGND VPWR VPWR _1833_/Y sky130_fd_sc_hd__xnor2_4
X_1764_ _1746_/A _1762_/Y _1763_/Y VGND VGND VPWR VPWR _1764_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_30_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1695_ _1696_/A _1695_/B VGND VGND VPWR VPWR _1695_/X sky130_fd_sc_hd__or2_4
X_2178_ _2181_/CLK _2178_/D VGND VGND VPWR VPWR _1609_/C sky130_fd_sc_hd__dfxtp_4
X_1129_ _1116_/C _1087_/Y _1091_/X _1090_/C _1126_/C VGND VGND VPWR VPWR _1129_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_25_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9_0_addressalyzerBlock.SPI_CLK clkbuf_4_9_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2225_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1480_ _1480_/A _1480_/B VGND VGND VPWR VPWR _1480_/X sky130_fd_sc_hd__and2_4
X_2101_ _2110_/CLK _1859_/Y VGND VGND VPWR VPWR _2101_/Q sky130_fd_sc_hd__dfxtp_4
X_2032_ _2027_/CLK _2032_/D VGND VGND VPWR VPWR HASH_ADDR[3] sky130_fd_sc_hd__dfxtp_4
X_1816_ _2121_/Q _1815_/X VGND VGND VPWR VPWR _1816_/X sky130_fd_sc_hd__xor2_4
X_1747_ _1739_/X _1930_/A _1746_/Y VGND VGND VPWR VPWR _1747_/Y sky130_fd_sc_hd__o21ai_4
X_1678_ _1963_/A _1678_/B VGND VGND VPWR VPWR _2162_/D sky130_fd_sc_hd__nor2_4
XFILLER_41_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1601_ _1600_/Y VGND VGND VPWR VPWR _1601_/Y sky130_fd_sc_hd__inv_2
X_1532_ _2198_/Q _1525_/X _1531_/X VGND VGND VPWR VPWR _1532_/X sky130_fd_sc_hd__o21a_4
X_1394_ _1313_/C _2117_/Q _1313_/B _1366_/A VGND VGND VPWR VPWR _1394_/X sky130_fd_sc_hd__a211o_4
X_1463_ _1387_/X _1463_/B VGND VGND VPWR VPWR _1463_/Y sky130_fd_sc_hd__nor2_4
X_2015_ _2016_/CLK _2015_/D VGND VGND VPWR VPWR _2015_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_23_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_m1_clk_local clkbuf_2_1_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_3_3_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_0_0_addressalyzerBlock.SPI_CLK clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_3_1_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
X_1515_ _1503_/X _1316_/A _1510_/X VGND VGND VPWR VPWR _1515_/X sky130_fd_sc_hd__o21a_4
XFILLER_55_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1377_ _1377_/A VGND VGND VPWR VPWR _1473_/B sky130_fd_sc_hd__buf_2
X_1446_ _1446_/A VGND VGND VPWR VPWR _1446_/X sky130_fd_sc_hd__buf_2
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1231_ _1159_/X _2065_/Q _1161_/X VGND VGND VPWR VPWR _1231_/Y sky130_fd_sc_hd__a21oi_4
X_1162_ _1159_/X _2066_/Q _1161_/X VGND VGND VPWR VPWR _1162_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_37_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1300_ _1298_/Y _1299_/Y _1339_/A VGND VGND VPWR VPWR _1300_/X sky130_fd_sc_hd__a21o_4
XFILLER_64_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1093_ _1058_/X _1076_/A _1091_/X _1090_/D _1092_/X VGND VGND VPWR VPWR _1093_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1995_ _2110_/CLK _1715_/A VGND VGND VPWR VPWR _2019_/D sky130_fd_sc_hd__dfxtp_4
X_1429_ _1427_/Y _1428_/X _1282_/C VGND VGND VPWR VPWR _1429_/X sky130_fd_sc_hd__o21a_4
XFILLER_28_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1780_ _1831_/A _1771_/Y _1838_/B VGND VGND VPWR VPWR _1825_/A sky130_fd_sc_hd__nor3_4
XFILLER_42_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1145_ _1145_/A VGND VGND VPWR VPWR _1377_/A sky130_fd_sc_hd__inv_2
XFILLER_37_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1214_ _1207_/C _1207_/D VGND VGND VPWR VPWR _1215_/B sky130_fd_sc_hd__nand2_4
XFILLER_1_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2194_ _2202_/CLK _1543_/X VGND VGND VPWR VPWR _2194_/Q sky130_fd_sc_hd__dfxtp_4
X_1076_ _1076_/A _1058_/X _1090_/B _1090_/D VGND VGND VPWR VPWR _1076_/X sky130_fd_sc_hd__and4_4
X_1978_ _1977_/Y M1_CLK_SELECT VGND VGND VPWR VPWR _1978_/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1832_ _2113_/Q _1843_/B _1836_/C _1831_/Y VGND VGND VPWR VPWR _1832_/Y sky130_fd_sc_hd__nand4_4
X_1901_ _1316_/Y _1885_/X _1888_/X _1351_/Y _1890_/X VGND VGND VPWR VPWR _1901_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_34_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1763_ _1763_/A _1757_/B _1763_/C VGND VGND VPWR VPWR _1763_/Y sky130_fd_sc_hd__nand3_4
X_1694_ _1038_/X VGND VGND VPWR VPWR _1696_/A sky130_fd_sc_hd__buf_2
X_2246_ _2013_/CLK _2246_/D VGND VGND VPWR VPWR _2246_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2177_ _2181_/CLK _2177_/D VGND VGND VPWR VPWR _1585_/B sky130_fd_sc_hd__dfxtp_4
X_1128_ _1128_/A _1128_/B VGND VGND VPWR VPWR _1128_/Y sky130_fd_sc_hd__nand2_4
X_1059_ _1090_/D _1484_/A _1058_/X _1105_/B VGND VGND VPWR VPWR _1060_/A sky130_fd_sc_hd__and4_4
Xclkbuf_4_14_0_addressalyzerBlock.SPI_CLK clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2243_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2100_ _2110_/CLK _1861_/Y VGND VGND VPWR VPWR _1857_/B sky130_fd_sc_hd__dfxtp_4
X_2031_ _2022_/CLK _2031_/D VGND VGND VPWR VPWR HASH_ADDR[2] sky130_fd_sc_hd__dfxtp_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1815_ _1825_/A _1813_/C _1813_/D VGND VGND VPWR VPWR _1815_/X sky130_fd_sc_hd__and3_4
XFILLER_15_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1746_ _1746_/A _1746_/B _1230_/A VGND VGND VPWR VPWR _1746_/Y sky130_fd_sc_hd__nand3_4
X_1677_ _1678_/B _1670_/B _1676_/Y VGND VGND VPWR VPWR _2163_/D sky130_fd_sc_hd__o21a_4
XFILLER_7_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2229_ _2243_/CLK _1252_/Y VGND VGND VPWR VPWR _1251_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_5_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1462_ _1462_/A VGND VGND VPWR VPWR _1463_/B sky130_fd_sc_hd__inv_2
X_1600_ _1600_/A _1599_/X _1596_/A VGND VGND VPWR VPWR _1600_/Y sky130_fd_sc_hd__nand3_4
X_1531_ _2199_/Q _1526_/X _1521_/X VGND VGND VPWR VPWR _1531_/X sky130_fd_sc_hd__o21a_4
X_1393_ _1391_/Y _1285_/X _1392_/Y VGND VGND VPWR VPWR _1393_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2014_ _2214_/CLK _1975_/X VGND VGND VPWR VPWR _1438_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1729_ _1914_/B _1728_/Y _1202_/Y _1265_/B _1365_/A VGND VGND VPWR VPWR _1729_/Y
+ sky130_fd_sc_hd__o41ai_4
XFILLER_58_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1445_ _1443_/X _1445_/B _1445_/C _1449_/C VGND VGND VPWR VPWR _1445_/Y sky130_fd_sc_hd__nand4_4
XFILLER_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1514_ _1573_/B _2198_/Q _1513_/X VGND VGND VPWR VPWR _1514_/X sky130_fd_sc_hd__o21a_4
XFILLER_55_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1376_ _1804_/C VGND VGND VPWR VPWR _1788_/A sky130_fd_sc_hd__inv_2
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1230_ _1230_/A _1230_/B VGND VGND VPWR VPWR _1230_/Y sky130_fd_sc_hd__nand2_4
X_1161_ _1161_/A VGND VGND VPWR VPWR _1161_/X sky130_fd_sc_hd__buf_2
XFILLER_1_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1092_ _1092_/A VGND VGND VPWR VPWR _1092_/X sky130_fd_sc_hd__buf_2
X_1994_ SCSN_fromHost VGND VGND VPWR VPWR SCSN_toClient sky130_fd_sc_hd__buf_2
XFILLER_20_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1428_ _1001_/A _1972_/C VGND VGND VPWR VPWR _1428_/X sky130_fd_sc_hd__or2_4
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1359_ _1359_/A _1358_/X VGND VGND VPWR VPWR _1359_/Y sky130_fd_sc_hd__nand2_4
XFILLER_43_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1213_ _1213_/A VGND VGND VPWR VPWR _1216_/A sky130_fd_sc_hd__inv_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1144_ _1311_/A _1144_/B VGND VGND VPWR VPWR _1145_/A sky130_fd_sc_hd__nor2_4
XFILLER_37_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2193_ _2013_/CLK _2193_/D VGND VGND VPWR VPWR _2193_/Q sky130_fd_sc_hd__dfxtp_4
X_1075_ _1105_/B VGND VGND VPWR VPWR _1090_/B sky130_fd_sc_hd__buf_2
X_1977_ M1_CLK_IN VGND VGND VPWR VPWR _1977_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1831_ _1831_/A VGND VGND VPWR VPWR _1831_/Y sky130_fd_sc_hd__inv_2
X_1900_ _1112_/Y _1898_/Y _1899_/Y VGND VGND VPWR VPWR _2087_/D sky130_fd_sc_hd__o21ai_4
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1762_ _1935_/B _1443_/X _1762_/C VGND VGND VPWR VPWR _1762_/Y sky130_fd_sc_hd__nand3_4
X_1693_ _1689_/A _1693_/B _1693_/C _1693_/D VGND VGND VPWR VPWR _1693_/X sky130_fd_sc_hd__and4_4
X_2176_ _2181_/CLK _2176_/D VGND VGND VPWR VPWR _1585_/A sky130_fd_sc_hd__dfxtp_4
X_2245_ _2243_/CLK _2245_/D VGND VGND VPWR VPWR _2245_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_15_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1127_ _2204_/Q _1123_/X _1126_/Y VGND VGND VPWR VPWR _1128_/A sky130_fd_sc_hd__a21o_4
X_1058_ _1058_/A VGND VGND VPWR VPWR _1058_/X sky130_fd_sc_hd__buf_2
XFILLER_31_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2030_ _2016_/CLK _2036_/Q VGND VGND VPWR VPWR HASH_ADDR[1] sky130_fd_sc_hd__dfxtp_4
XFILLER_47_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1814_ _1814_/A _1813_/Y VGND VGND VPWR VPWR _2122_/D sky130_fd_sc_hd__xnor2_4
XFILLER_30_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1745_ _1633_/A _1740_/X _1892_/A VGND VGND VPWR VPWR _1930_/A sky130_fd_sc_hd__nand3_4
X_1676_ _1678_/B _1670_/B _1101_/X VGND VGND VPWR VPWR _1676_/Y sky130_fd_sc_hd__a21oi_4
X_2228_ _2050_/CLK _2228_/D VGND VGND VPWR VPWR _1274_/B sky130_fd_sc_hd__dfxtp_4
X_2159_ _2153_/CLK _2159_/D VGND VGND VPWR VPWR _2159_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_0_0_addressalyzerBlock.SPI_CLK clkbuf_3_1_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_4_1_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_13_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1392_ _1180_/B _2045_/Q _1188_/X VGND VGND VPWR VPWR _1392_/Y sky130_fd_sc_hd__o21ai_4
X_1461_ _1459_/Y _1460_/Y _1723_/A VGND VGND VPWR VPWR _1461_/X sky130_fd_sc_hd__a21o_4
X_1530_ _2199_/Q _1525_/X _1529_/X VGND VGND VPWR VPWR _2200_/D sky130_fd_sc_hd__o21a_4
XFILLER_8_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2013_ _2013_/CLK _1957_/Y VGND VGND VPWR VPWR _1451_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_50_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1728_ _1845_/A VGND VGND VPWR VPWR _1728_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1659_ _1659_/A VGND VGND VPWR VPWR _2168_/D sky130_fd_sc_hd__inv_2
XFILLER_41_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1375_ _1343_/X _1373_/Y _1374_/Y VGND VGND VPWR VPWR _1375_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_4_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1513_ _1503_/X _1753_/C _1510_/X VGND VGND VPWR VPWR _1513_/X sky130_fd_sc_hd__o21a_4
X_1444_ _1451_/B VGND VGND VPWR VPWR _1445_/C sky130_fd_sc_hd__inv_2
XFILLER_23_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1160_ _1175_/A VGND VGND VPWR VPWR _1161_/A sky130_fd_sc_hd__inv_2
X_1091_ _1090_/B VGND VGND VPWR VPWR _1091_/X sky130_fd_sc_hd__buf_2
XFILLER_60_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1993_ SCLK_fromHost VGND VGND VPWR VPWR SCLK_toClient sky130_fd_sc_hd__buf_2
XFILLER_13_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1358_ _1757_/C _1230_/B _1161_/X _1357_/Y VGND VGND VPWR VPWR _1358_/X sky130_fd_sc_hd__a211o_4
X_1427_ _1436_/A _2007_/Q VGND VGND VPWR VPWR _1427_/Y sky130_fd_sc_hd__nor2_4
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1289_ _1084_/A _1104_/Y _1288_/X VGND VGND VPWR VPWR _1289_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_46_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1212_ _1829_/B VGND VGND VPWR VPWR _1849_/A sky130_fd_sc_hd__inv_2
X_2192_ _2013_/CLK _1552_/Y VGND VGND VPWR VPWR _1545_/B sky130_fd_sc_hd__dfxtp_4
X_1143_ _2220_/Q VGND VGND VPWR VPWR _1144_/B sky130_fd_sc_hd__inv_2
XFILLER_37_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1074_ _1069_/Y _1073_/Y _1040_/X VGND VGND VPWR VPWR _2238_/D sky130_fd_sc_hd__a21oi_4
XFILLER_18_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1976_ EXT_RESET_N_fromHost VGND VGND VPWR VPWR _2003_/D sky130_fd_sc_hd__inv_2
XFILLER_29_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1830_ _1829_/X VGND VGND VPWR VPWR _1843_/B sky130_fd_sc_hd__buf_2
XFILLER_30_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1761_ _1746_/A _1759_/Y _1760_/Y VGND VGND VPWR VPWR _2133_/D sky130_fd_sc_hd__o21ai_4
X_1692_ _1692_/A VGND VGND VPWR VPWR _1693_/C sky130_fd_sc_hd__inv_2
X_1126_ _1126_/A _1482_/B _1126_/C _1125_/Y VGND VGND VPWR VPWR _1126_/Y sky130_fd_sc_hd__nor4_4
X_2175_ _2181_/CLK _1635_/Y VGND VGND VPWR VPWR _1577_/A sky130_fd_sc_hd__dfxtp_4
X_2244_ _2243_/CLK _2244_/D VGND VGND VPWR VPWR _2244_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_33_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1057_ _1057_/A _1057_/B _1057_/C _1124_/A VGND VGND VPWR VPWR _1090_/D sky130_fd_sc_hd__and4_4
XFILLER_21_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1959_ _1696_/A _1036_/B _1972_/C _1971_/C _1958_/Y VGND VGND VPWR VPWR _2007_/D
+ sky130_fd_sc_hd__o41ai_4
XFILLER_56_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_6_0_m1_clk_local clkbuf_2_3_0_m1_clk_local/X VGND VGND VPWR VPWR _2127_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1813_ _2121_/Q _1827_/B _1813_/C _1813_/D VGND VGND VPWR VPWR _1813_/Y sky130_fd_sc_hd__nand4_4
X_1744_ _1739_/X _1928_/A _1743_/Y VGND VGND VPWR VPWR _1744_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_30_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1675_ _1674_/X _1307_/B _1675_/C VGND VGND VPWR VPWR _2164_/D sky130_fd_sc_hd__and3_4
X_2089_ _2042_/CLK _1893_/Y VGND VGND VPWR VPWR _2089_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2227_ _2214_/CLK _1287_/Y VGND VGND VPWR VPWR _1147_/A sky130_fd_sc_hd__dfxtp_4
X_2158_ _2216_/CLK _1685_/X VGND VGND VPWR VPWR _2158_/Q sky130_fd_sc_hd__dfxtp_4
X_1109_ _1120_/A _1106_/X _1126_/A _1116_/C VGND VGND VPWR VPWR _1109_/Y sky130_fd_sc_hd__nand4_4
XFILLER_53_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1391_ _1386_/X _1390_/X VGND VGND VPWR VPWR _1391_/Y sky130_fd_sc_hd__nand2_4
X_1460_ _1460_/A _1355_/X VGND VGND VPWR VPWR _1460_/Y sky130_fd_sc_hd__nand2_4
XFILLER_4_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2012_ _2013_/CLK _1965_/Y VGND VGND VPWR VPWR _1964_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_35_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1727_ _1313_/C _1827_/A _1313_/B _1198_/A VGND VGND VPWR VPWR _1727_/X sky130_fd_sc_hd__a211o_4
X_1658_ _1648_/X _1647_/Y _1657_/Y VGND VGND VPWR VPWR _1659_/A sky130_fd_sc_hd__o21ai_4
X_1589_ _2181_/Q _1600_/A _1589_/C _1596_/C VGND VGND VPWR VPWR _1589_/Y sky130_fd_sc_hd__nand4_4
XFILLER_41_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1512_ _1573_/B _2199_/Q _1511_/X VGND VGND VPWR VPWR _1512_/X sky130_fd_sc_hd__o21a_4
X_1374_ _1274_/A _2219_/Q VGND VGND VPWR VPWR _1374_/Y sky130_fd_sc_hd__nand2_4
X_1443_ _1927_/D VGND VGND VPWR VPWR _1443_/X sky130_fd_sc_hd__buf_2
XFILLER_48_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1090_ _1087_/Y _1090_/B _1090_/C _1090_/D VGND VGND VPWR VPWR _1090_/X sky130_fd_sc_hd__and4_4
X_1992_ MOSI_fromHost VGND VGND VPWR VPWR MOSI_toClient sky130_fd_sc_hd__buf_2
X_1357_ _1355_/X _1357_/B VGND VGND VPWR VPWR _1357_/Y sky130_fd_sc_hd__nor2_4
XFILLER_28_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1288_ _1087_/A _1104_/A _1086_/X _1049_/X _1298_/C VGND VGND VPWR VPWR _1288_/X
+ sky130_fd_sc_hd__o41a_4
X_1426_ _2216_/Q VGND VGND VPWR VPWR _1426_/Y sky130_fd_sc_hd__inv_2
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1211_ _1211_/A VGND VGND VPWR VPWR _1829_/B sky130_fd_sc_hd__buf_2
X_2191_ _2013_/CLK _2191_/D VGND VGND VPWR VPWR _1545_/C sky130_fd_sc_hd__dfxtp_4
X_1142_ _1138_/Y _1140_/Y _1141_/Y VGND VGND VPWR VPWR _1142_/Y sky130_fd_sc_hd__a21oi_4
X_1073_ _1070_/X _1072_/Y _1969_/B VGND VGND VPWR VPWR _1073_/Y sky130_fd_sc_hd__o21ai_4
X_1975_ _1974_/X _1436_/Y _1701_/A VGND VGND VPWR VPWR _1975_/X sky130_fd_sc_hd__o21a_4
X_1409_ _1407_/Y _1233_/X _1408_/Y VGND VGND VPWR VPWR _1409_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_0_0_addressalyzerBlock.SPI_CLK clkbuf_4_1_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2207_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_42_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1760_ _1763_/A _1757_/B _2133_/Q VGND VGND VPWR VPWR _1760_/Y sky130_fd_sc_hd__nand3_4
X_1691_ _1957_/A _1692_/A _1693_/D _1693_/B VGND VGND VPWR VPWR _1691_/Y sky130_fd_sc_hd__nor4_4
X_2243_ _2243_/CLK _1019_/Y VGND VGND VPWR VPWR _2243_/Q sky130_fd_sc_hd__dfxtp_4
X_2174_ _2181_/CLK _1638_/Y VGND VGND VPWR VPWR _1576_/A sky130_fd_sc_hd__dfxtp_4
X_1125_ _1090_/B _1104_/Y _1088_/X _1084_/A VGND VGND VPWR VPWR _1125_/Y sky130_fd_sc_hd__nand4_4
X_1056_ _1092_/A VGND VGND VPWR VPWR _1056_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1889_ _1897_/C _1218_/X _1195_/X _1927_/D _1292_/X VGND VGND VPWR VPWR _1889_/X
+ sky130_fd_sc_hd__a41o_4
X_1958_ _1753_/A _1061_/A _1001_/A _1325_/X VGND VGND VPWR VPWR _1958_/Y sky130_fd_sc_hd__nand4_4
XFILLER_56_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_5_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1812_ _1825_/A VGND VGND VPWR VPWR _1827_/B sky130_fd_sc_hd__buf_2
X_1743_ _1746_/A _1746_/B _1156_/A VGND VGND VPWR VPWR _1743_/Y sky130_fd_sc_hd__nand3_4
XFILLER_7_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1674_ _2162_/Q _1670_/B _2164_/Q VGND VGND VPWR VPWR _1674_/X sky130_fd_sc_hd__a21o_4
X_2226_ _2214_/CLK _1295_/Y VGND VGND VPWR VPWR _1147_/B sky130_fd_sc_hd__dfxtp_4
X_2088_ _2083_/CLK _2088_/D VGND VGND VPWR VPWR _1258_/A sky130_fd_sc_hd__dfxtp_4
X_2157_ _2153_/CLK _2157_/D VGND VGND VPWR VPWR _2157_/Q sky130_fd_sc_hd__dfxtp_4
X_1039_ _1038_/X VGND VGND VPWR VPWR _1039_/X sky130_fd_sc_hd__buf_2
X_1108_ _1124_/A VGND VGND VPWR VPWR _1116_/C sky130_fd_sc_hd__buf_2
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1390_ _2133_/Q _1230_/B _1161_/A _1389_/Y VGND VGND VPWR VPWR _1390_/X sky130_fd_sc_hd__a211o_4
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2011_ _2214_/CLK _1968_/X VGND VGND VPWR VPWR _1451_/C sky130_fd_sc_hd__dfxtp_4
X_1726_ _2115_/Q VGND VGND VPWR VPWR _1827_/A sky130_fd_sc_hd__buf_2
X_1657_ _1647_/Y _1648_/X _1293_/X VGND VGND VPWR VPWR _1657_/Y sky130_fd_sc_hd__a21oi_4
X_1588_ _1574_/Y _1588_/B VGND VGND VPWR VPWR _1600_/A sky130_fd_sc_hd__nor2_4
X_2209_ _2207_/CLK _1506_/X VGND VGND VPWR VPWR _1741_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1442_ _1737_/D VGND VGND VPWR VPWR _1927_/D sky130_fd_sc_hd__buf_2
X_1511_ _1503_/X _1894_/A _1510_/X VGND VGND VPWR VPWR _1511_/X sky130_fd_sc_hd__o21a_4
XFILLER_4_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1373_ THREAD_COUNT[3] _1345_/X _1369_/Y _1372_/Y VGND VGND VPWR VPWR _1373_/Y sky130_fd_sc_hd__a22oi_4
X_1709_ _1217_/X _1708_/A _1215_/Y _1708_/X VGND VGND VPWR VPWR _1709_/X sky130_fd_sc_hd__a211o_4
XFILLER_54_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1991_ EXT_RESET_N_fromHost VGND VGND VPWR VPWR EXT_RESET_N_toClient sky130_fd_sc_hd__buf_2
X_1425_ _1343_/X _1423_/Y _1424_/Y VGND VGND VPWR VPWR _2217_/D sky130_fd_sc_hd__o21ai_4
XFILLER_55_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1287_ _1277_/Y _1284_/Y _1286_/X VGND VGND VPWR VPWR _1287_/Y sky130_fd_sc_hd__a21oi_4
X_1356_ _1356_/A VGND VGND VPWR VPWR _1357_/B sky130_fd_sc_hd__inv_2
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2190_ _2016_/CLK _2190_/D VGND VGND VPWR VPWR _1981_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_49_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1210_ _1203_/Y _1833_/A _1209_/X VGND VGND VPWR VPWR _1210_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_37_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1072_ _1076_/A _1061_/D _1126_/C VGND VGND VPWR VPWR _1072_/Y sky130_fd_sc_hd__a21oi_4
X_1141_ _1091_/X _1128_/B _1031_/X VGND VGND VPWR VPWR _1141_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_18_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1974_ _1436_/A _1451_/A _1451_/C VGND VGND VPWR VPWR _1974_/X sky130_fd_sc_hd__o21a_4
XFILLER_56_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1408_ _1171_/X _2036_/D _1172_/X VGND VGND VPWR VPWR _1408_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_45_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1339_ _1339_/A _1144_/B VGND VGND VPWR VPWR _1339_/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1690_ _1957_/A _2146_/Q _1689_/B VGND VGND VPWR VPWR _1690_/Y sky130_fd_sc_hd__nor3_4
X_2242_ _2243_/CLK _1023_/Y VGND VGND VPWR VPWR _2242_/Q sky130_fd_sc_hd__dfxtp_4
X_2173_ _2173_/CLK _1640_/Y VGND VGND VPWR VPWR _2173_/Q sky130_fd_sc_hd__dfxtp_4
X_1055_ _1054_/Y VGND VGND VPWR VPWR _1092_/A sky130_fd_sc_hd__buf_2
XFILLER_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1124_ _1124_/A VGND VGND VPWR VPWR _1482_/B sky130_fd_sc_hd__inv_2
X_1957_ _1957_/A _1445_/B _1092_/X VGND VGND VPWR VPWR _1957_/Y sky130_fd_sc_hd__nor3_4
XFILLER_21_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1888_ _1905_/A VGND VGND VPWR VPWR _1888_/X sky130_fd_sc_hd__buf_2
XFILLER_0_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1811_ _1803_/A _1787_/Y VGND VGND VPWR VPWR _2123_/D sky130_fd_sc_hd__xor2_4
XFILLER_30_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1742_ _1739_/A VGND VGND VPWR VPWR _1746_/A sky130_fd_sc_hd__buf_2
X_1673_ _1581_/D _1671_/Y _1672_/Y VGND VGND VPWR VPWR _1673_/X sky130_fd_sc_hd__o21a_4
X_2225_ _2225_/CLK _2225_/D VGND VGND VPWR VPWR _1149_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_53_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2087_ _2069_/CLK _2087_/D VGND VGND VPWR VPWR _1999_/D sky130_fd_sc_hd__dfxtp_4
X_1038_ _1886_/A VGND VGND VPWR VPWR _1038_/X sky130_fd_sc_hd__buf_2
X_2156_ _2153_/CLK _2156_/D VGND VGND VPWR VPWR _1456_/B sky130_fd_sc_hd__dfxtp_4
X_1107_ _1057_/C VGND VGND VPWR VPWR _1126_/A sky130_fd_sc_hd__buf_2
XFILLER_21_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2010_ _2225_/CLK _2010_/D VGND VGND VPWR VPWR _1278_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_50_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_2_0_m1_clk_local clkbuf_3_3_0_m1_clk_local/A VGND VGND VPWR VPWR _2022_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1725_ _1711_/Y _1723_/Y _1724_/Y VGND VGND VPWR VPWR _1725_/Y sky130_fd_sc_hd__o21ai_4
X_1587_ _1609_/C _1584_/Y _1587_/C _1609_/D VGND VGND VPWR VPWR _1588_/B sky130_fd_sc_hd__nand4_4
X_1656_ _1957_/A _1656_/B _1655_/Y VGND VGND VPWR VPWR _2169_/D sky130_fd_sc_hd__nor3_4
X_2139_ _2077_/CLK _1736_/Y VGND VGND VPWR VPWR _2139_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_26_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2208_ _2207_/CLK _2208_/D VGND VGND VPWR VPWR _1892_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1441_ _1436_/Y _1438_/Y _1440_/X VGND VGND VPWR VPWR _1441_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1510_ _1633_/A VGND VGND VPWR VPWR _1510_/X sky130_fd_sc_hd__buf_2
XFILLER_63_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1372_ _1209_/X _1856_/A _1345_/X VGND VGND VPWR VPWR _1372_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_31_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1708_ _1708_/A THREAD_COUNT[0] _1708_/C VGND VGND VPWR VPWR _1708_/X sky130_fd_sc_hd__and3_4
XFILLER_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1639_ _1607_/X _1646_/C _1031_/X VGND VGND VPWR VPWR _1639_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1990_ _1988_/Y _1964_/A _1989_/Y VGND VGND VPWR VPWR _2246_/D sky130_fd_sc_hd__a21oi_4
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1355_ _1405_/A VGND VGND VPWR VPWR _1355_/X sky130_fd_sc_hd__buf_2
X_1424_ _1480_/A _1424_/B VGND VGND VPWR VPWR _1424_/Y sky130_fd_sc_hd__nand2_4
XFILLER_63_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1286_ _1283_/X _1285_/X _1446_/A VGND VGND VPWR VPWR _1286_/X sky130_fd_sc_hd__a21o_4
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_5_0_addressalyzerBlock.SPI_CLK clkbuf_3_2_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2042_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_37_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1140_ _1907_/A _1123_/X _1079_/X VGND VGND VPWR VPWR _1140_/Y sky130_fd_sc_hd__a21oi_4
X_1071_ _1092_/A VGND VGND VPWR VPWR _1126_/C sky130_fd_sc_hd__buf_2
XFILLER_18_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1973_ _1553_/Y _2005_/Q _1696_/A _1972_/X VGND VGND VPWR VPWR _2005_/D sky130_fd_sc_hd__a211o_4
X_1407_ _2084_/Q VGND VGND VPWR VPWR _1407_/Y sky130_fd_sc_hd__inv_2
X_1338_ _1907_/A _1279_/Y _1337_/X _1283_/A VGND VGND VPWR VPWR _1338_/X sky130_fd_sc_hd__a211o_4
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1269_ _1203_/Y _1839_/A _1209_/X VGND VGND VPWR VPWR _1269_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_36_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2241_ _2243_/CLK _1027_/Y VGND VGND VPWR VPWR _1024_/A sky130_fd_sc_hd__dfxtp_4
X_2172_ _2173_/CLK _1646_/X VGND VGND VPWR VPWR _2172_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1123_ _1278_/B VGND VGND VPWR VPWR _1123_/X sky130_fd_sc_hd__buf_2
X_1054_ _1449_/A _1309_/A VGND VGND VPWR VPWR _1054_/Y sky130_fd_sc_hd__nor2_4
X_1887_ _1886_/Y VGND VGND VPWR VPWR _1905_/A sky130_fd_sc_hd__inv_2
X_1956_ _1720_/B _1948_/X _1907_/A _1943_/A VGND VGND VPWR VPWR _2059_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1810_ _2124_/Q _1804_/B VGND VGND VPWR VPWR _1810_/X sky130_fd_sc_hd__xor2_4
X_1741_ _1917_/A _1740_/X _1741_/C VGND VGND VPWR VPWR _1928_/A sky130_fd_sc_hd__nand3_4
X_1672_ _1678_/B _1670_/B _2164_/Q _1581_/D _1039_/X VGND VGND VPWR VPWR _1672_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_7_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2224_ _2214_/CLK _2224_/D VGND VGND VPWR VPWR _1149_/B sky130_fd_sc_hd__dfxtp_4
X_2155_ _2013_/CLK _1690_/Y VGND VGND VPWR VPWR _1972_/C sky130_fd_sc_hd__dfxtp_4
X_1106_ _1106_/A VGND VGND VPWR VPWR _1106_/X sky130_fd_sc_hd__buf_2
X_2086_ _2042_/CLK _1901_/Y VGND VGND VPWR VPWR _2086_/Q sky130_fd_sc_hd__dfxtp_4
X_1037_ _2004_/Q VGND VGND VPWR VPWR _1886_/A sky130_fd_sc_hd__buf_2
X_1939_ _1904_/Y _1934_/Y _1732_/X _1404_/Y _1935_/Y VGND VGND VPWR VPWR _2068_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_44_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0_addressalyzerBlock.SPI_CLK clkbuf_0_addressalyzerBlock.SPI_CLK/X VGND
+ VGND VPWR VPWR clkbuf_2_3_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_35_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1724_ _1187_/A _1769_/A _1153_/Y VGND VGND VPWR VPWR _1724_/Y sky130_fd_sc_hd__a21oi_4
X_1655_ _1647_/Y _1648_/X _1643_/X VGND VGND VPWR VPWR _1655_/Y sky130_fd_sc_hd__a21oi_4
X_1586_ _1585_/Y VGND VGND VPWR VPWR _1609_/D sky130_fd_sc_hd__inv_2
X_2069_ _2069_/CLK _1938_/Y VGND VGND VPWR VPWR _1380_/A sky130_fd_sc_hd__dfxtp_4
X_2138_ _2083_/CLK _1744_/Y VGND VGND VPWR VPWR _1156_/A sky130_fd_sc_hd__dfxtp_4
X_2207_ _2207_/CLK _1512_/X VGND VGND VPWR VPWR _1748_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_5_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1371_ _1370_/Y VGND VGND VPWR VPWR _1856_/A sky130_fd_sc_hd__buf_2
X_1440_ _1886_/C _1298_/C _1496_/B _1451_/A VGND VGND VPWR VPWR _1440_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1707_ _1342_/A VGND VGND VPWR VPWR _2140_/D sky130_fd_sc_hd__inv_2
X_1638_ _1638_/A VGND VGND VPWR VPWR _1638_/Y sky130_fd_sc_hd__inv_2
X_1569_ _2186_/Q _2187_/Q VGND VGND VPWR VPWR _1569_/X sky130_fd_sc_hd__or2_4
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1354_ _1350_/X _1353_/Y _1175_/X VGND VGND VPWR VPWR _1359_/A sky130_fd_sc_hd__a21o_4
X_1285_ _1263_/B VGND VGND VPWR VPWR _1285_/X sky130_fd_sc_hd__buf_2
X_1423_ THREAD_COUNT[1] _1345_/X _1420_/Y _1422_/X VGND VGND VPWR VPWR _1423_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_51_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_10_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2153_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1070_ _1067_/Y VGND VGND VPWR VPWR _1070_/X sky130_fd_sc_hd__buf_2
X_1972_ _1971_/Y _1004_/A _1972_/C VGND VGND VPWR VPWR _1972_/X sky130_fd_sc_hd__and3_4
X_1406_ _2076_/Q _1154_/X _1166_/X _1405_/Y VGND VGND VPWR VPWR _1406_/X sky130_fd_sc_hd__a211o_4
X_1268_ _1153_/Y _1266_/Y _1267_/X VGND VGND VPWR VPWR _1268_/Y sky130_fd_sc_hd__o21ai_4
X_1337_ _1449_/A _1309_/A _1144_/B VGND VGND VPWR VPWR _1337_/X sky130_fd_sc_hd__o21a_4
XFILLER_61_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1199_ _1195_/X _1814_/A _1196_/X _1473_/C VGND VGND VPWR VPWR _1199_/X sky130_fd_sc_hd__a211o_4
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2171_ _2173_/CLK _2171_/D VGND VGND VPWR VPWR _1583_/C sky130_fd_sc_hd__dfxtp_4
X_1122_ _1118_/Y _1119_/Y _1121_/X VGND VGND VPWR VPWR _2234_/D sky130_fd_sc_hd__a21oi_4
X_2240_ _2243_/CLK _1033_/Y VGND VGND VPWR VPWR _2240_/Q sky130_fd_sc_hd__dfxtp_4
X_1053_ _1052_/X VGND VGND VPWR VPWR _1076_/A sky130_fd_sc_hd__buf_2
X_1886_ _1886_/A _1886_/B _1886_/C VGND VGND VPWR VPWR _1886_/Y sky130_fd_sc_hd__nor3_4
X_1955_ _1412_/B _1949_/X _1762_/C _1950_/X VGND VGND VPWR VPWR _2060_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1740_ _1927_/D VGND VGND VPWR VPWR _1740_/X sky130_fd_sc_hd__buf_2
XFILLER_30_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1671_ _1675_/C VGND VGND VPWR VPWR _1671_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2085_ _2083_/CLK _1903_/Y VGND VGND VPWR VPWR _2085_/Q sky130_fd_sc_hd__dfxtp_4
X_2223_ _2077_/CLK _1324_/Y VGND VGND VPWR VPWR _1048_/A sky130_fd_sc_hd__dfxtp_4
X_1105_ _1104_/Y _1105_/B _1147_/A _1147_/B VGND VGND VPWR VPWR _1106_/A sky130_fd_sc_hd__and4_4
X_2154_ _2202_/CLK _1691_/Y VGND VGND VPWR VPWR _1526_/A sky130_fd_sc_hd__dfxtp_4
X_1036_ _2139_/Q _1036_/B VGND VGND VPWR VPWR _1036_/Y sky130_fd_sc_hd__nand2_4
X_1938_ _1902_/Y _1934_/Y _1732_/X _1380_/Y _1935_/Y VGND VGND VPWR VPWR _1938_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1869_ _1867_/A _1867_/B _2097_/Q VGND VGND VPWR VPWR _1869_/Y sky130_fd_sc_hd__nand3_4
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1723_ _1723_/A _1722_/Y VGND VGND VPWR VPWR _1723_/Y sky130_fd_sc_hd__nor2_4
X_1654_ _1654_/A VGND VGND VPWR VPWR _1957_/A sky130_fd_sc_hd__buf_2
X_1585_ _1585_/A _1585_/B VGND VGND VPWR VPWR _1585_/Y sky130_fd_sc_hd__nand2_4
X_2206_ _2202_/CLK _1514_/X VGND VGND VPWR VPWR _1753_/C sky130_fd_sc_hd__dfxtp_4
X_2068_ _2056_/CLK _2068_/D VGND VGND VPWR VPWR _1404_/A sky130_fd_sc_hd__dfxtp_4
X_2137_ _2137_/CLK _1747_/Y VGND VGND VPWR VPWR _1230_/A sky130_fd_sc_hd__dfxtp_4
X_1019_ _1017_/Y _1003_/X _1018_/Y VGND VGND VPWR VPWR _1019_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_1_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1370_ _2102_/Q VGND VGND VPWR VPWR _1370_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1706_ _1318_/X _1323_/C _1333_/Y _1334_/Y _1335_/X VGND VGND VPWR VPWR _1706_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1637_ _1621_/B _1619_/Y _1636_/Y VGND VGND VPWR VPWR _1638_/A sky130_fd_sc_hd__o21ai_4
X_1568_ _1570_/A SPI_CLK_RESET_N _1562_/Y _1568_/D VGND VGND VPWR VPWR _2188_/D sky130_fd_sc_hd__and4_4
XFILLER_39_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1499_ _1426_/Y _1499_/B VGND VGND VPWR VPWR _1499_/Y sky130_fd_sc_hd__nand2_4
XFILLER_54_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1422_ _1857_/B _1365_/A _1421_/Y VGND VGND VPWR VPWR _1422_/X sky130_fd_sc_hd__o21a_4
XFILLER_9_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1353_ _1351_/Y _1233_/X _1352_/Y VGND VGND VPWR VPWR _1353_/Y sky130_fd_sc_hd__o21ai_4
X_1284_ _1741_/C _1279_/Y _1283_/X VGND VGND VPWR VPWR _1284_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_36_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0999_ _2244_/Q _1034_/A _0998_/X VGND VGND VPWR VPWR _0999_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1971_ _1971_/A _1320_/Y _1971_/C VGND VGND VPWR VPWR _1971_/Y sky130_fd_sc_hd__nand3_4
X_1405_ _1405_/A _1404_/Y VGND VGND VPWR VPWR _1405_/Y sky130_fd_sc_hd__nor2_4
X_1198_ _1198_/A VGND VGND VPWR VPWR _1473_/C sky130_fd_sc_hd__buf_2
X_1267_ _1195_/X _1783_/A _1196_/X _1473_/C VGND VGND VPWR VPWR _1267_/X sky130_fd_sc_hd__a211o_4
X_1336_ _1318_/X _1323_/C _1333_/Y _1334_/Y _1335_/X VGND VGND VPWR VPWR _1336_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_51_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_addressalyzerBlock.SPI_CLK _1982_/Y VGND VGND VPWR VPWR clkbuf_0_addressalyzerBlock.SPI_CLK/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_19_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2170_ _2173_/CLK _2170_/D VGND VGND VPWR VPWR _1644_/A sky130_fd_sc_hd__dfxtp_4
X_1121_ _1070_/X _1120_/Y _1446_/A VGND VGND VPWR VPWR _1121_/X sky130_fd_sc_hd__a21o_4
X_1052_ _1050_/Y _1723_/A _1147_/B _1149_/A VGND VGND VPWR VPWR _1052_/X sky130_fd_sc_hd__and4_4
XFILLER_33_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1954_ _1389_/B _1949_/X _1902_/A _1950_/X VGND VGND VPWR VPWR _1954_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_2_1_0_addressalyzerBlock.SPI_CLK clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_3_2_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
X_1885_ _1473_/B VGND VGND VPWR VPWR _1885_/X sky130_fd_sc_hd__buf_2
XFILLER_56_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1319_ _1449_/A VGND VGND VPWR VPWR _1971_/A sky130_fd_sc_hd__inv_2
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1670_ _1678_/B _1670_/B _2164_/Q VGND VGND VPWR VPWR _1675_/C sky130_fd_sc_hd__nand3_4
XFILLER_7_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2222_ _2069_/CLK _1332_/Y VGND VGND VPWR VPWR _1184_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2084_ _2042_/CLK _1906_/Y VGND VGND VPWR VPWR _2084_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1104_ _1104_/A _1086_/A _1048_/Y VGND VGND VPWR VPWR _1104_/Y sky130_fd_sc_hd__nor3_4
X_2153_ _2153_/CLK _1693_/X VGND VGND VPWR VPWR _1011_/A sky130_fd_sc_hd__dfxtp_4
X_1035_ _1001_/A VGND VGND VPWR VPWR _1036_/B sky130_fd_sc_hd__buf_2
XFILLER_61_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1937_ _1316_/Y _1934_/Y _1732_/X _1348_/Y _1935_/Y VGND VGND VPWR VPWR _2070_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1799_ _1799_/A _1799_/B VGND VGND VPWR VPWR _1799_/Y sky130_fd_sc_hd__nand2_4
X_1868_ _1928_/A _1865_/X _1867_/Y VGND VGND VPWR VPWR _1868_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_44_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1722_ _1718_/Y _1161_/X _1721_/X VGND VGND VPWR VPWR _1722_/Y sky130_fd_sc_hd__a21boi_4
X_1584_ _1575_/Y _1608_/B _1577_/Y _1583_/Y VGND VGND VPWR VPWR _1584_/Y sky130_fd_sc_hd__nor4_4
X_1653_ _1644_/X _1656_/B _1652_/Y VGND VGND VPWR VPWR _2170_/D sky130_fd_sc_hd__o21a_4
X_2205_ _2202_/CLK _2205_/D VGND VGND VPWR VPWR _1316_/A sky130_fd_sc_hd__dfxtp_4
X_2136_ _2142_/CLK _1752_/Y VGND VGND VPWR VPWR _1253_/A sky130_fd_sc_hd__dfxtp_4
X_2067_ _2137_/CLK _1941_/X VGND VGND VPWR VPWR _2067_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_34_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1018_ _1480_/B _1004_/X _1008_/X VGND VGND VPWR VPWR _1018_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_19_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1705_ _1318_/X _1323_/C _1327_/Y _1328_/Y _1331_/X VGND VGND VPWR VPWR _2142_/D
+ sky130_fd_sc_hd__a41oi_4
XFILLER_31_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1567_ _2186_/Q _2187_/Q _1562_/C VGND VGND VPWR VPWR _1568_/D sky130_fd_sc_hd__a21o_4
XFILLER_58_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1636_ _1619_/Y _1621_/B _1293_/X VGND VGND VPWR VPWR _1636_/Y sky130_fd_sc_hd__a21oi_4
X_2119_ _2127_/CLK _2119_/D VGND VGND VPWR VPWR _1817_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_54_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1498_ _2216_/Q _1498_/B _2144_/Q _1493_/X VGND VGND VPWR VPWR _1498_/Y sky130_fd_sc_hd__nand4_4
XFILLER_13_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_15_0_addressalyzerBlock.SPI_CLK clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2050_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_57_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1421_ _1345_/X VGND VGND VPWR VPWR _1421_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1352_ _1164_/X _2094_/Q _1172_/X VGND VGND VPWR VPWR _1352_/Y sky130_fd_sc_hd__a21oi_4
X_1283_ _1283_/A VGND VGND VPWR VPWR _1283_/X sky130_fd_sc_hd__buf_2
XFILLER_36_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0998_ _2245_/Q _0997_/X VGND VGND VPWR VPWR _0998_/X sky130_fd_sc_hd__or2_4
X_1619_ _1607_/X _1646_/C VGND VGND VPWR VPWR _1619_/Y sky130_fd_sc_hd__nor2_4
XFILLER_54_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1970_ _1971_/A _1960_/X _1969_/Y VGND VGND VPWR VPWR _2008_/D sky130_fd_sc_hd__o21ai_4
XFILLER_18_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1404_ _1404_/A VGND VGND VPWR VPWR _1404_/Y sky130_fd_sc_hd__inv_2
X_1335_ _1339_/A _1218_/X _1654_/A VGND VGND VPWR VPWR _1335_/X sky130_fd_sc_hd__a21o_4
XFILLER_56_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1266_ _1264_/Y _1188_/X _1265_/Y VGND VGND VPWR VPWR _1266_/Y sky130_fd_sc_hd__a21oi_4
X_1197_ _1153_/B VGND VGND VPWR VPWR _1198_/A sky130_fd_sc_hd__buf_2
XFILLER_36_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1051_ _1147_/A VGND VGND VPWR VPWR _1723_/A sky130_fd_sc_hd__buf_2
XFILLER_18_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1120_ _1120_/A VGND VGND VPWR VPWR _1120_/Y sky130_fd_sc_hd__inv_2
X_1884_ _1940_/A _1867_/A _1883_/Y VGND VGND VPWR VPWR _1884_/Y sky130_fd_sc_hd__o21ai_4
X_1953_ _1357_/B _1949_/X _1316_/A _1950_/X VGND VGND VPWR VPWR _2062_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1318_ _1318_/A VGND VGND VPWR VPWR _1318_/X sky130_fd_sc_hd__buf_2
XFILLER_64_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1249_ _1248_/Y _1209_/A _1272_/B VGND VGND VPWR VPWR _1249_/X sky130_fd_sc_hd__a21o_4
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2221_ _2077_/CLK _1336_/Y VGND VGND VPWR VPWR _1205_/A sky130_fd_sc_hd__dfxtp_4
X_2152_ _2153_/CLK _1695_/X VGND VGND VPWR VPWR _1692_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2083_ _2083_/CLK _2083_/D VGND VGND VPWR VPWR _1715_/A sky130_fd_sc_hd__dfxtp_4
X_1103_ _1057_/B VGND VGND VPWR VPWR _1120_/A sky130_fd_sc_hd__buf_2
X_1034_ _1034_/A _1004_/X _1028_/A VGND VGND VPWR VPWR _1034_/Y sky130_fd_sc_hd__nand3_4
XFILLER_21_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1936_ _1112_/Y _1934_/Y _1732_/X _1463_/B _1935_/Y VGND VGND VPWR VPWR _1936_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1867_ _1867_/A _1867_/B _2098_/Q VGND VGND VPWR VPWR _1867_/Y sky130_fd_sc_hd__nand3_4
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1798_ _1809_/B _1789_/X _1804_/C _1791_/Y _2129_/Q VGND VGND VPWR VPWR _1799_/A
+ sky130_fd_sc_hd__a41o_4
XFILLER_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1721_ _2131_/Q _1387_/X _1161_/A _1720_/Y VGND VGND VPWR VPWR _1721_/X sky130_fd_sc_hd__a211o_4
XFILLER_11_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1652_ _1648_/X _1647_/Y _1643_/X _1644_/X _1039_/X VGND VGND VPWR VPWR _1652_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1583_ _1644_/A _1656_/B _1583_/C _2172_/Q VGND VGND VPWR VPWR _1583_/Y sky130_fd_sc_hd__nand4_4
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2135_ _2142_/CLK _2135_/D VGND VGND VPWR VPWR _1460_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_26_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2204_ _2202_/CLK _1518_/X VGND VGND VPWR VPWR _2204_/Q sky130_fd_sc_hd__dfxtp_4
X_2066_ _2069_/CLK _1945_/Y VGND VGND VPWR VPWR _2066_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_41_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1017_ _2242_/Q _1034_/A _1016_/X VGND VGND VPWR VPWR _1017_/Y sky130_fd_sc_hd__o21ai_4
X_1919_ _1112_/Y _1918_/A _1918_/Y VGND VGND VPWR VPWR _1919_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_1_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1704_ _1689_/A ID_fromClient VGND VGND VPWR VPWR _2143_/D sky130_fd_sc_hd__and2_4
X_1566_ _1566_/A SPI_CLK_RESET_N _1570_/A VGND VGND VPWR VPWR _1566_/X sky130_fd_sc_hd__and3_4
X_1635_ _1577_/Y _1632_/Y _1634_/Y VGND VGND VPWR VPWR _1635_/Y sky130_fd_sc_hd__a21oi_4
X_1497_ _1495_/Y _1496_/Y _1446_/X VGND VGND VPWR VPWR _2211_/D sky130_fd_sc_hd__a21oi_4
XFILLER_54_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2118_ _2121_/CLK _2118_/D VGND VGND VPWR VPWR _1781_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_39_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2049_ _2137_/CLK _2057_/Q VGND VGND VPWR VPWR _2049_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1351_ _2086_/Q VGND VGND VPWR VPWR _1351_/Y sky130_fd_sc_hd__inv_2
X_1420_ _1420_/A _1397_/B _1420_/C VGND VGND VPWR VPWR _1420_/Y sky130_fd_sc_hd__nand3_4
XFILLER_63_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1282_ _1282_/A _1318_/A _1282_/C VGND VGND VPWR VPWR _1283_/A sky130_fd_sc_hd__nand3_4
X_1618_ _1583_/Y VGND VGND VPWR VPWR _1646_/C sky130_fd_sc_hd__buf_2
X_0997_ _1011_/A VGND VGND VPWR VPWR _0997_/X sky130_fd_sc_hd__buf_2
XFILLER_39_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1549_ _1549_/A VGND VGND VPWR VPWR _1549_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_1_0_addressalyzerBlock.SPI_CLK clkbuf_3_1_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_4_3_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_40_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1265_ _1802_/A _1265_/B _1732_/A VGND VGND VPWR VPWR _1265_/Y sky130_fd_sc_hd__nor3_4
X_1403_ _1402_/Y _1189_/A _1191_/A _1377_/A _1366_/A VGND VGND VPWR VPWR _1403_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1334_ _1217_/X _1708_/C _1298_/C VGND VGND VPWR VPWR _1334_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_51_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1196_ _1311_/A VGND VGND VPWR VPWR _1196_/X sky130_fd_sc_hd__buf_2
XFILLER_59_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_0_m1_clk_local clkbuf_2_1_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_3_1_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1050_ _1086_/A _1049_/X VGND VGND VPWR VPWR _1050_/Y sky130_fd_sc_hd__nor2_4
XFILLER_33_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1952_ _1487_/Y _1949_/X _1753_/C _1950_/X VGND VGND VPWR VPWR _2063_/D sky130_fd_sc_hd__a2bb2o_4
X_1883_ _1864_/Y _1899_/B _1883_/C VGND VGND VPWR VPWR _1883_/Y sky130_fd_sc_hd__nand3_4
XFILLER_56_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1248_ _1829_/C VGND VGND VPWR VPWR _1248_/Y sky130_fd_sc_hd__inv_2
X_1317_ _1215_/A _1126_/C _1313_/Y _1316_/Y _1279_/A VGND VGND VPWR VPWR _1317_/Y
+ sky130_fd_sc_hd__o32ai_4
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1179_ _1263_/B VGND VGND VPWR VPWR _1180_/B sky130_fd_sc_hd__buf_2
XFILLER_12_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2082_ _2083_/CLK _2082_/D VGND VGND VPWR VPWR _2082_/Q sky130_fd_sc_hd__dfxtp_4
X_2220_ _2077_/CLK _1342_/Y VGND VGND VPWR VPWR _2220_/Q sky130_fd_sc_hd__dfxtp_4
X_2151_ _2225_/CLK _2151_/D VGND VGND VPWR VPWR _1695_/B sky130_fd_sc_hd__dfxtp_4
X_1102_ _1101_/X VGND VGND VPWR VPWR _1963_/A sky130_fd_sc_hd__buf_2
XFILLER_46_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1033_ _1029_/Y _1964_/A _1032_/Y VGND VGND VPWR VPWR _1033_/Y sky130_fd_sc_hd__a21oi_4
X_1797_ _1402_/Y _1803_/A _1787_/Y VGND VGND VPWR VPWR _1809_/B sky130_fd_sc_hd__nor3_4
X_1935_ _1935_/A _1935_/B VGND VGND VPWR VPWR _1935_/Y sky130_fd_sc_hd__nand2_4
X_1866_ _1864_/Y VGND VGND VPWR VPWR _1867_/A sky130_fd_sc_hd__buf_2
XFILLER_52_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1720_ _1154_/X _1720_/B VGND VGND VPWR VPWR _1720_/Y sky130_fd_sc_hd__nor2_4
X_1651_ _1583_/C _1649_/X _1650_/Y VGND VGND VPWR VPWR _2171_/D sky130_fd_sc_hd__o21a_4
X_1582_ _1582_/A _1582_/B _1647_/A _1582_/D VGND VGND VPWR VPWR _1656_/B sky130_fd_sc_hd__nor4_4
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2065_ _2069_/CLK _1947_/Y VGND VGND VPWR VPWR _2065_/Q sky130_fd_sc_hd__dfxtp_4
X_2134_ _2142_/CLK _2134_/D VGND VGND VPWR VPWR _1757_/C sky130_fd_sc_hd__dfxtp_4
X_2203_ _2202_/CLK _1520_/X VGND VGND VPWR VPWR _1904_/A sky130_fd_sc_hd__dfxtp_4
X_1016_ _2243_/Q _1016_/B VGND VGND VPWR VPWR _1016_/X sky130_fd_sc_hd__or2_4
X_1849_ _1849_/A _1779_/B VGND VGND VPWR VPWR _1850_/A sky130_fd_sc_hd__xor2_4
X_1918_ _1918_/A _1918_/B _1918_/C VGND VGND VPWR VPWR _1918_/Y sky130_fd_sc_hd__nand3_4
XFILLER_57_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1703_ _1689_/A _2143_/Q VGND VGND VPWR VPWR _1703_/X sky130_fd_sc_hd__and2_4
X_1634_ _1607_/X _1608_/B _1577_/Y _1646_/C _1753_/A VGND VGND VPWR VPWR _1634_/Y
+ sky130_fd_sc_hd__o41ai_4
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1565_ _1565_/A VGND VGND VPWR VPWR _1570_/A sky130_fd_sc_hd__inv_2
X_1496_ _1426_/Y _1496_/B VGND VGND VPWR VPWR _1496_/Y sky130_fd_sc_hd__nand2_4
X_2048_ _2056_/CLK _2048_/D VGND VGND VPWR VPWR _1263_/A sky130_fd_sc_hd__dfxtp_4
X_2117_ _2121_/CLK _1824_/Y VGND VGND VPWR VPWR _2117_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1350_ HASH_LED _1154_/X _1166_/X _1349_/Y VGND VGND VPWR VPWR _1350_/X sky130_fd_sc_hd__a211o_4
X_1281_ _1281_/A VGND VGND VPWR VPWR _1282_/C sky130_fd_sc_hd__inv_2
XFILLER_63_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0996_ _0996_/A VGND VGND VPWR VPWR _1034_/A sky130_fd_sc_hd__buf_2
X_1617_ _1616_/X _1307_/B _1595_/C VGND VGND VPWR VPWR _2179_/D sky130_fd_sc_hd__and3_4
X_1479_ _1474_/X _1476_/Y _1478_/Y VGND VGND VPWR VPWR _1479_/X sky130_fd_sc_hd__a21o_4
X_1548_ _1011_/A _1545_/C VGND VGND VPWR VPWR _1549_/A sky130_fd_sc_hd__nand2_4
XFILLER_54_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1402_ _2124_/Q VGND VGND VPWR VPWR _1402_/Y sky130_fd_sc_hd__inv_2
X_1264_ _1088_/X _1262_/Y _1263_/X VGND VGND VPWR VPWR _1264_/Y sky130_fd_sc_hd__o21ai_4
X_1333_ _1325_/X _1123_/X _1762_/C VGND VGND VPWR VPWR _1333_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_51_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1195_ _1312_/A VGND VGND VPWR VPWR _1195_/X sky130_fd_sc_hd__buf_2
XFILLER_24_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1882_ _1762_/Y _1867_/A _1881_/Y VGND VGND VPWR VPWR _2092_/D sky130_fd_sc_hd__o21ai_4
X_1951_ _1490_/Y _1949_/X _1894_/A _1950_/X VGND VGND VPWR VPWR _2064_/D sky130_fd_sc_hd__a2bb2o_4
X_1247_ _1203_/Y _2113_/Q _1209_/X VGND VGND VPWR VPWR _1247_/Y sky130_fd_sc_hd__a21oi_4
X_1178_ _1147_/A VGND VGND VPWR VPWR _1263_/B sky130_fd_sc_hd__inv_2
X_1316_ _1316_/A VGND VGND VPWR VPWR _1316_/Y sky130_fd_sc_hd__inv_2
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2081_ _2042_/CLK _1912_/Y VGND VGND VPWR VPWR _1232_/A sky130_fd_sc_hd__dfxtp_4
X_2150_ _2153_/CLK _2150_/D VGND VGND VPWR VPWR _1682_/B sky130_fd_sc_hd__dfxtp_4
X_1101_ _1038_/X VGND VGND VPWR VPWR _1101_/X sky130_fd_sc_hd__buf_2
X_1032_ _1424_/B _1003_/A _1031_/X VGND VGND VPWR VPWR _1032_/Y sky130_fd_sc_hd__o21ai_4
X_1934_ _1934_/A VGND VGND VPWR VPWR _1934_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1796_ _1796_/A _1796_/B VGND VGND VPWR VPWR _1796_/Y sky130_fd_sc_hd__nor2_4
X_1865_ _1864_/Y VGND VGND VPWR VPWR _1865_/X sky130_fd_sc_hd__buf_2
XFILLER_44_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1650_ _1643_/X _1642_/Y _1644_/X _1583_/C _1039_/X VGND VGND VPWR VPWR _1650_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1581_ _2162_/Q _1581_/B _2164_/Q _1581_/D VGND VGND VPWR VPWR _1582_/D sky130_fd_sc_hd__nand4_4
XFILLER_7_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2202_ _2202_/CLK _1523_/X VGND VGND VPWR VPWR _1139_/A sky130_fd_sc_hd__dfxtp_4
X_2133_ _2142_/CLK _2133_/D VGND VGND VPWR VPWR _2133_/Q sky130_fd_sc_hd__dfxtp_4
X_2064_ _2142_/CLK _2064_/D VGND VGND VPWR VPWR _1490_/A sky130_fd_sc_hd__dfxtp_4
X_1015_ _1013_/Y _1003_/X _1014_/Y VGND VGND VPWR VPWR _2244_/D sky130_fd_sc_hd__a21oi_4
X_1917_ _1917_/A VGND VGND VPWR VPWR _1918_/B sky130_fd_sc_hd__buf_2
X_1779_ _1211_/A _1779_/B _1836_/B _1836_/C VGND VGND VPWR VPWR _1838_/B sky130_fd_sc_hd__nand4_4
X_1848_ _1847_/X VGND VGND VPWR VPWR _1848_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_1_0_addressalyzerBlock.SPI_CLK clkbuf_4_1_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2137_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1564_ _1562_/Y _1563_/A _1563_/Y VGND VGND VPWR VPWR _1566_/A sky130_fd_sc_hd__a21o_4
X_1633_ _1633_/A VGND VGND VPWR VPWR _1753_/A sky130_fd_sc_hd__buf_2
X_1702_ _1701_/A _1693_/C VGND VGND VPWR VPWR _1702_/Y sky130_fd_sc_hd__nand2_4
XFILLER_39_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1495_ _1495_/A _2216_/Q _2144_/Q VGND VGND VPWR VPWR _1495_/Y sky130_fd_sc_hd__nand3_4
X_2116_ _2121_/CLK _1826_/X VGND VGND VPWR VPWR _2116_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_54_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2047_ _2216_/CLK _2055_/Q VGND VGND VPWR VPWR _2047_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_addressalyzerBlock.SPI_CLK clkbuf_2_3_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1280_ _1280_/A _1066_/A VGND VGND VPWR VPWR _1281_/A sky130_fd_sc_hd__nor2_4
XFILLER_51_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0995_ _1011_/A VGND VGND VPWR VPWR _0996_/A sky130_fd_sc_hd__inv_2
XFILLER_59_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1616_ _1609_/A _1621_/C _1609_/C _1609_/D _1587_/C VGND VGND VPWR VPWR _1616_/X
+ sky130_fd_sc_hd__a41o_4
X_1547_ _1544_/Y _1545_/Y _1546_/Y VGND VGND VPWR VPWR _2193_/D sky130_fd_sc_hd__a21oi_4
XFILLER_54_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1478_ _1477_/Y _1397_/B _1222_/Y VGND VGND VPWR VPWR _1478_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_39_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1401_ _1343_/X _1399_/Y _1400_/Y VGND VGND VPWR VPWR _2218_/D sky130_fd_sc_hd__o21ai_4
X_1263_ _1263_/A _1263_/B VGND VGND VPWR VPWR _1263_/X sky130_fd_sc_hd__or2_4
X_1194_ _2220_/Q VGND VGND VPWR VPWR _1312_/A sky130_fd_sc_hd__buf_2
X_1332_ _1318_/X _1323_/C _1327_/Y _1328_/Y _1331_/X VGND VGND VPWR VPWR _1332_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_17_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1950_ _1943_/A VGND VGND VPWR VPWR _1950_/X sky130_fd_sc_hd__buf_2
XFILLER_33_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1881_ _1874_/A _1899_/B _2036_/D VGND VGND VPWR VPWR _1881_/Y sky130_fd_sc_hd__nand3_4
X_1315_ _1314_/X _1283_/X _1215_/A VGND VGND VPWR VPWR _1315_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_56_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1246_ _1153_/Y _1244_/Y _1245_/X VGND VGND VPWR VPWR _1246_/Y sky130_fd_sc_hd__o21ai_4
X_1177_ _1156_/Y _1162_/Y _1176_/Y VGND VGND VPWR VPWR _1177_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2080_ _2042_/CLK _1913_/Y VGND VGND VPWR VPWR ID_toHost sky130_fd_sc_hd__dfxtp_4
XFILLER_53_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1100_ _1094_/Y _1096_/Y _1099_/X VGND VGND VPWR VPWR _2236_/D sky130_fd_sc_hd__a21oi_4
X_1031_ _1750_/A VGND VGND VPWR VPWR _1031_/X sky130_fd_sc_hd__buf_2
XFILLER_61_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1933_ _1935_/A _1341_/C _2072_/Q _1185_/A _1932_/Y VGND VGND VPWR VPWR _1933_/X
+ sky130_fd_sc_hd__a32o_4
X_1795_ _1795_/A _1799_/B VGND VGND VPWR VPWR _1796_/B sky130_fd_sc_hd__nor2_4
X_1864_ _1864_/A VGND VGND VPWR VPWR _1864_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1229_ _1229_/A _1229_/B VGND VGND VPWR VPWR _1229_/Y sky130_fd_sc_hd__nand2_4
XFILLER_32_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1580_ _1660_/A _1580_/B VGND VGND VPWR VPWR _1647_/A sky130_fd_sc_hd__nand2_4
X_2132_ _2142_/CLK _1764_/Y VGND VGND VPWR VPWR _1763_/C sky130_fd_sc_hd__dfxtp_4
X_2201_ _2207_/CLK _1528_/X VGND VGND VPWR VPWR _2201_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_34_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2063_ _2142_/CLK _2063_/D VGND VGND VPWR VPWR _1487_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1014_ _1274_/B _1004_/X _1008_/X VGND VGND VPWR VPWR _1014_/Y sky130_fd_sc_hd__o21ai_4
X_1847_ _1728_/Y _1836_/A VGND VGND VPWR VPWR _1847_/X sky130_fd_sc_hd__xor2_4
X_1916_ _1924_/A VGND VGND VPWR VPWR _1918_/A sky130_fd_sc_hd__buf_2
X_1778_ _1777_/Y VGND VGND VPWR VPWR _1836_/C sky130_fd_sc_hd__inv_2
XFILLER_57_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1701_ _1701_/A _1689_/B VGND VGND VPWR VPWR _1701_/Y sky130_fd_sc_hd__nand2_4
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1563_ _1563_/A _1570_/C VGND VGND VPWR VPWR _1563_/Y sky130_fd_sc_hd__nor2_4
X_1632_ _1609_/A VGND VGND VPWR VPWR _1632_/Y sky130_fd_sc_hd__inv_2
X_1494_ _1498_/B _1493_/X _1061_/D VGND VGND VPWR VPWR _1495_/A sky130_fd_sc_hd__a21o_4
X_2115_ _2121_/CLK _1827_/X VGND VGND VPWR VPWR _2115_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_54_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2046_ _2216_/CLK _2054_/Q VGND VGND VPWR VPWR _2046_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_5_0_m1_clk_local clkbuf_3_4_0_m1_clk_local/A VGND VGND VPWR VPWR _2027_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1477_ _2103_/Q VGND VGND VPWR VPWR _1477_/Y sky130_fd_sc_hd__inv_2
X_1615_ _1577_/A VGND VGND VPWR VPWR _1621_/C sky130_fd_sc_hd__buf_2
X_1546_ _1546_/A _1457_/A VGND VGND VPWR VPWR _1546_/Y sky130_fd_sc_hd__nand2_4
XFILLER_39_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2029_ _2027_/CLK _2029_/D VGND VGND VPWR VPWR HASH_ADDR[0] sky130_fd_sc_hd__dfxtp_4
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1331_ _1339_/A _1897_/C _1654_/A VGND VGND VPWR VPWR _1331_/X sky130_fd_sc_hd__a21o_4
X_1400_ _1274_/A _1400_/B VGND VGND VPWR VPWR _1400_/Y sky130_fd_sc_hd__nand2_4
X_1193_ _1181_/Y _1188_/X _1192_/Y VGND VGND VPWR VPWR _1193_/Y sky130_fd_sc_hd__a21oi_4
X_1262_ _1253_/Y _1254_/Y _1261_/Y VGND VGND VPWR VPWR _1262_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_36_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1529_ _2200_/Q _1526_/X _1521_/X VGND VGND VPWR VPWR _1529_/X sky130_fd_sc_hd__o21a_4
XFILLER_19_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1880_ _1759_/Y _1867_/A _1879_/Y VGND VGND VPWR VPWR _2093_/D sky130_fd_sc_hd__o21ai_4
XFILLER_14_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1314_ _1436_/A _1451_/A _1313_/Y VGND VGND VPWR VPWR _1314_/X sky130_fd_sc_hd__o21a_4
XFILLER_52_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1245_ _1195_/X _2121_/Q _1196_/X _1473_/C VGND VGND VPWR VPWR _1245_/X sky130_fd_sc_hd__a211o_4
X_1176_ _1168_/Y _1174_/Y _1175_/X VGND VGND VPWR VPWR _1176_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_20_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1030_ _1004_/A VGND VGND VPWR VPWR _1964_/A sky130_fd_sc_hd__buf_2
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1932_ _1932_/A VGND VGND VPWR VPWR _1932_/Y sky130_fd_sc_hd__inv_2
X_1863_ _1419_/C _1863_/B _1152_/D _1737_/D VGND VGND VPWR VPWR _1864_/A sky130_fd_sc_hd__and4_4
XFILLER_14_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1794_ _2129_/Q _1788_/Y _1789_/X _1791_/Y VGND VGND VPWR VPWR _1799_/B sky130_fd_sc_hd__nand4_4
XFILLER_37_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1228_ _1274_/A _2230_/Q VGND VGND VPWR VPWR _1229_/B sky130_fd_sc_hd__nand2_4
X_1159_ _1170_/A VGND VGND VPWR VPWR _1159_/X sky130_fd_sc_hd__buf_2
XFILLER_20_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2131_ _2137_/CLK _1768_/Y VGND VGND VPWR VPWR _2131_/Q sky130_fd_sc_hd__dfxtp_4
X_2062_ _2142_/CLK _2062_/D VGND VGND VPWR VPWR _1356_/A sky130_fd_sc_hd__dfxtp_4
X_2200_ _2207_/CLK _2200_/D VGND VGND VPWR VPWR _2200_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_4_6_0_addressalyzerBlock.SPI_CLK clkbuf_4_7_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2069_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_34_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1013_ _2243_/Q _1034_/A _1012_/X VGND VGND VPWR VPWR _1013_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_19_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1777_ _1842_/A _2109_/Q VGND VGND VPWR VPWR _1777_/Y sky130_fd_sc_hd__nand2_4
X_1846_ _2108_/Q _1846_/B VGND VGND VPWR VPWR _1846_/Y sky130_fd_sc_hd__xnor2_4
X_1915_ _1914_/Y VGND VGND VPWR VPWR _1924_/A sky130_fd_sc_hd__inv_2
XFILLER_57_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1700_ _1689_/A MOSI_fromHost VGND VGND VPWR VPWR _2147_/D sky130_fd_sc_hd__and2_4
X_1631_ _1585_/A _1584_/Y _1630_/Y VGND VGND VPWR VPWR _2176_/D sky130_fd_sc_hd__o21a_4
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1562_ _2186_/Q _2187_/Q _1562_/C VGND VGND VPWR VPWR _1562_/Y sky130_fd_sc_hd__nand3_4
X_1493_ _1488_/X _1489_/Y _1491_/Y _1493_/D VGND VGND VPWR VPWR _1493_/X sky130_fd_sc_hd__and4_4
X_2045_ _2056_/CLK _2053_/Q VGND VGND VPWR VPWR _2045_/Q sky130_fd_sc_hd__dfxtp_4
X_2114_ _2121_/CLK _1833_/Y VGND VGND VPWR VPWR _1833_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_62_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1829_ _1851_/B _1829_/B _1829_/C _1836_/B VGND VGND VPWR VPWR _1829_/X sky130_fd_sc_hd__and4_4
XFILLER_57_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1614_ _1574_/Y _1595_/C _1613_/Y VGND VGND VPWR VPWR _1614_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_8_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1476_ _1203_/Y _1838_/A _1209_/A VGND VGND VPWR VPWR _1476_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_39_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1545_ _0997_/X _1545_/B _1545_/C VGND VGND VPWR VPWR _1545_/Y sky130_fd_sc_hd__nand3_4
XFILLER_54_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2028_ _2110_/CLK _2067_/Q VGND VGND VPWR VPWR _2027_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1261_ _1257_/Y _1260_/Y _1175_/X VGND VGND VPWR VPWR _1261_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_30_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1330_ _1292_/X VGND VGND VPWR VPWR _1654_/A sky130_fd_sc_hd__buf_2
X_1192_ _2130_/Q _1265_/B _1732_/A VGND VGND VPWR VPWR _1192_/Y sky130_fd_sc_hd__nor3_4
XFILLER_36_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1459_ _1159_/X _1487_/A _1161_/A VGND VGND VPWR VPWR _1459_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1528_ _2200_/Q _1525_/X _1527_/X VGND VGND VPWR VPWR _1528_/X sky130_fd_sc_hd__o21a_4
XFILLER_42_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1244_ _1242_/Y _1188_/X _1243_/Y VGND VGND VPWR VPWR _1244_/Y sky130_fd_sc_hd__a21oi_4
X_1313_ _1886_/B _1313_/B _1313_/C VGND VGND VPWR VPWR _1313_/Y sky130_fd_sc_hd__nand3_4
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1175_ _1175_/A VGND VGND VPWR VPWR _1175_/X sky130_fd_sc_hd__buf_2
XFILLER_24_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1793_ _2130_/Q VGND VGND VPWR VPWR _1795_/A sky130_fd_sc_hd__inv_2
X_1931_ _1935_/A _1341_/C _2073_/Q _1185_/A _1930_/Y VGND VGND VPWR VPWR _1931_/X
+ sky130_fd_sc_hd__a32o_4
X_1862_ _1922_/C _1857_/C VGND VGND VPWR VPWR _2099_/D sky130_fd_sc_hd__xor2_4
XFILLER_6_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1158_ _1171_/A VGND VGND VPWR VPWR _1170_/A sky130_fd_sc_hd__buf_2
X_1227_ _1480_/A VGND VGND VPWR VPWR _1274_/A sky130_fd_sc_hd__buf_2
XFILLER_40_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1089_ _1088_/X VGND VGND VPWR VPWR _1090_/C sky130_fd_sc_hd__buf_2
XFILLER_20_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_11_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2013_/CLK sky130_fd_sc_hd__clkbuf_1
X_2130_ _2127_/CLK _1796_/Y VGND VGND VPWR VPWR _2130_/Q sky130_fd_sc_hd__dfxtp_4
X_2061_ _2142_/CLK _1954_/X VGND VGND VPWR VPWR _1388_/A sky130_fd_sc_hd__dfxtp_4
X_1012_ _2244_/Q _1016_/B VGND VGND VPWR VPWR _1012_/X sky130_fd_sc_hd__or2_4
X_1914_ _1886_/A _1914_/B _1886_/C _1909_/X VGND VGND VPWR VPWR _1914_/Y sky130_fd_sc_hd__nor4_4
XFILLER_22_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1845_ _1845_/A _1851_/B _1829_/B _1829_/C VGND VGND VPWR VPWR _1846_/B sky130_fd_sc_hd__nand4_4
X_1776_ _1776_/A VGND VGND VPWR VPWR _1836_/B sky130_fd_sc_hd__inv_2
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1630_ _1621_/B _1619_/Y _1621_/C _1585_/A _1039_/X VGND VGND VPWR VPWR _1630_/Y
+ sky130_fd_sc_hd__a41oi_4
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1561_ _1560_/X VGND VGND VPWR VPWR _2190_/D sky130_fd_sc_hd__inv_2
X_1492_ _1482_/B _2060_/Q _1057_/C _1389_/B VGND VGND VPWR VPWR _1493_/D sky130_fd_sc_hd__a22oi_4
X_2113_ _2121_/CLK _1837_/Y VGND VGND VPWR VPWR _2113_/Q sky130_fd_sc_hd__dfxtp_4
X_2044_ _2083_/CLK _2044_/D VGND VGND VPWR VPWR _2044_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_62_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1828_ _1856_/A _1774_/C _1856_/B VGND VGND VPWR VPWR _1851_/B sky130_fd_sc_hd__nor3_4
X_1759_ _1935_/B _1443_/X _1902_/A VGND VGND VPWR VPWR _1759_/Y sky130_fd_sc_hd__nand3_4
XFILLER_1_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1613_ _1574_/Y _1595_/C _1031_/X VGND VGND VPWR VPWR _1613_/Y sky130_fd_sc_hd__o21ai_4
X_1544_ _2193_/Q VGND VGND VPWR VPWR _1544_/Y sky130_fd_sc_hd__inv_2
X_1475_ _1770_/B VGND VGND VPWR VPWR _1838_/A sky130_fd_sc_hd__inv_2
XFILLER_39_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2027_ _2027_/CLK _2027_/D VGND VGND VPWR VPWR MACRO_RD_SELECT sky130_fd_sc_hd__dfxtp_4
XFILLER_49_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1191_ _1191_/A VGND VGND VPWR VPWR _1732_/A sky130_fd_sc_hd__buf_2
X_1260_ _1258_/Y _1170_/X _1259_/Y VGND VGND VPWR VPWR _1260_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_51_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_1_0_m1_clk_local clkbuf_3_1_0_m1_clk_local/A VGND VGND VPWR VPWR _2173_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1527_ _2201_/Q _1526_/X _1521_/X VGND VGND VPWR VPWR _1527_/X sky130_fd_sc_hd__o21a_4
X_1389_ _1387_/X _1389_/B VGND VGND VPWR VPWR _1389_/Y sky130_fd_sc_hd__nor2_4
X_1458_ _1546_/A _1458_/B VGND VGND VPWR VPWR _2213_/D sky130_fd_sc_hd__nor2_4
XFILLER_42_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1243_ _2129_/Q _1265_/B _1732_/A VGND VGND VPWR VPWR _1243_/Y sky130_fd_sc_hd__nor3_4
X_1174_ _1169_/Y _1170_/X _1173_/Y VGND VGND VPWR VPWR _1174_/Y sky130_fd_sc_hd__o21ai_4
X_1312_ _1312_/A VGND VGND VPWR VPWR _1313_/C sky130_fd_sc_hd__buf_2
XFILLER_2_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1930_ _1930_/A VGND VGND VPWR VPWR _1930_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1792_ _2129_/Q _1788_/Y _1789_/X _1791_/Y _2130_/Q VGND VGND VPWR VPWR _1796_/A
+ sky130_fd_sc_hd__a41oi_4
X_1861_ _1857_/B _1861_/B VGND VGND VPWR VPWR _1861_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_6_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1157_ _1347_/A VGND VGND VPWR VPWR _1171_/A sky130_fd_sc_hd__inv_2
XFILLER_37_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1226_ _1216_/A VGND VGND VPWR VPWR _1480_/A sky130_fd_sc_hd__buf_2
XFILLER_52_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1088_ _1723_/A VGND VGND VPWR VPWR _1088_/X sky130_fd_sc_hd__buf_2
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2060_ _2142_/CLK _2060_/D VGND VGND VPWR VPWR _2060_/Q sky130_fd_sc_hd__dfxtp_4
X_1011_ _1011_/A VGND VGND VPWR VPWR _1016_/B sky130_fd_sc_hd__buf_2
XFILLER_19_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1913_ _1894_/Y _1909_/X _1905_/X _1255_/Y _1910_/X VGND VGND VPWR VPWR _1913_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1844_ _1844_/A VGND VGND VPWR VPWR _1844_/Y sky130_fd_sc_hd__inv_2
X_1775_ _2108_/Q _1845_/A VGND VGND VPWR VPWR _1776_/A sky130_fd_sc_hd__nand2_4
XFILLER_8_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2189_ _2016_/CLK _1566_/X VGND VGND VPWR VPWR _1563_/A sky130_fd_sc_hd__dfxtp_4
X_1209_ _1209_/A VGND VGND VPWR VPWR _1209_/X sky130_fd_sc_hd__buf_2
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1560_ _1981_/A _1565_/A _1559_/Y VGND VGND VPWR VPWR _1560_/X sky130_fd_sc_hd__a21o_4
X_2112_ _2121_/CLK _2112_/D VGND VGND VPWR VPWR _1839_/A sky130_fd_sc_hd__dfxtp_4
X_1491_ _1120_/Y _1356_/A _1058_/X _1490_/Y VGND VGND VPWR VPWR _1491_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_3_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2043_ _2042_/CLK _2043_/D VGND VGND VPWR VPWR _2043_/Q sky130_fd_sc_hd__dfxtp_4
X_1827_ _1827_/A _1827_/B VGND VGND VPWR VPWR _1827_/X sky130_fd_sc_hd__xor2_4
X_1758_ _1739_/X _1756_/Y _1757_/Y VGND VGND VPWR VPWR _2134_/D sky130_fd_sc_hd__o21ai_4
X_1689_ _1689_/A _1689_/B _2146_/Q VGND VGND VPWR VPWR _2156_/D sky130_fd_sc_hd__and3_4
XFILLER_57_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_0_addressalyzerBlock.SPI_CLK clkbuf_2_3_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_48_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1474_ _1470_/Y _1471_/X _1203_/Y _1473_/Y VGND VGND VPWR VPWR _1474_/X sky130_fd_sc_hd__a211o_4
X_1543_ _1525_/A _2148_/Q _1542_/X VGND VGND VPWR VPWR _1543_/X sky130_fd_sc_hd__o21a_4
X_1612_ _1612_/A VGND VGND VPWR VPWR _1612_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2026_ _2022_/CLK _2026_/D VGND VGND VPWR VPWR DATA_TO_HASH[7] sky130_fd_sc_hd__dfxtp_4
XFILLER_35_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1190_ _1186_/B VGND VGND VPWR VPWR _1191_/A sky130_fd_sc_hd__buf_2
X_1457_ _1457_/A VGND VGND VPWR VPWR _1458_/B sky130_fd_sc_hd__inv_2
X_1526_ _1526_/A VGND VGND VPWR VPWR _1526_/X sky130_fd_sc_hd__buf_2
X_1388_ _1388_/A VGND VGND VPWR VPWR _1389_/B sky130_fd_sc_hd__inv_2
XFILLER_27_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2009_ _2225_/CLK _2009_/D VGND VGND VPWR VPWR _1325_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_46_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1311_ _1311_/A VGND VGND VPWR VPWR _1313_/B sky130_fd_sc_hd__buf_2
XFILLER_64_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1242_ _1088_/X _1240_/Y _1241_/X VGND VGND VPWR VPWR _1242_/Y sky130_fd_sc_hd__o21ai_4
X_1173_ _1171_/X _2098_/Q _1172_/X VGND VGND VPWR VPWR _1173_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_2_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1509_ _1863_/B VGND VGND VPWR VPWR _1633_/A sky130_fd_sc_hd__buf_2
XFILLER_46_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1860_ _1922_/C _1857_/C VGND VGND VPWR VPWR _1861_/B sky130_fd_sc_hd__nand2_4
X_1791_ _1790_/Y VGND VGND VPWR VPWR _1791_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1225_ _1200_/Y _1210_/Y _1224_/X VGND VGND VPWR VPWR _1229_/A sky130_fd_sc_hd__a21o_4
X_1156_ _1156_/A _1230_/B VGND VGND VPWR VPWR _1156_/Y sky130_fd_sc_hd__nand2_4
XFILLER_37_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1087_ _1087_/A _1104_/A _1086_/X _1049_/X VGND VGND VPWR VPWR _1087_/Y sky130_fd_sc_hd__nor4_4
X_1989_ _2230_/Q _1003_/A _1746_/B VGND VGND VPWR VPWR _1989_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1010_ _0999_/Y _1003_/X _1009_/Y VGND VGND VPWR VPWR _2245_/D sky130_fd_sc_hd__a21oi_4
X_1843_ _2109_/Q _1843_/B VGND VGND VPWR VPWR _1844_/A sky130_fd_sc_hd__xnor2_4
X_1912_ _1892_/Y _1909_/X _1905_/X _1232_/Y _1910_/X VGND VGND VPWR VPWR _1912_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_8_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1774_ _1248_/Y _1370_/Y _1774_/C _1856_/B VGND VGND VPWR VPWR _1779_/B sky130_fd_sc_hd__nor4_4
X_1208_ _1207_/X VGND VGND VPWR VPWR _1209_/A sky130_fd_sc_hd__buf_2
X_2188_ _2016_/CLK _2188_/D VGND VGND VPWR VPWR _1562_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_25_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1139_ _1139_/A VGND VGND VPWR VPWR _1907_/A sky130_fd_sc_hd__buf_2
XFILLER_56_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1490_ _1490_/A VGND VGND VPWR VPWR _1490_/Y sky130_fd_sc_hd__inv_2
X_2042_ _2042_/CLK DATA_AVAILABLE VGND VGND VPWR VPWR _2042_/Q sky130_fd_sc_hd__dfxtp_4
X_2111_ _2121_/CLK _2111_/D VGND VGND VPWR VPWR _1770_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_39_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1826_ _2116_/Q _1825_/X VGND VGND VPWR VPWR _1826_/X sky130_fd_sc_hd__xor2_4
XFILLER_30_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1757_ _1763_/A _1757_/B _1757_/C VGND VGND VPWR VPWR _1757_/Y sky130_fd_sc_hd__nand3_4
X_1688_ _2145_/Q VGND VGND VPWR VPWR _1689_/B sky130_fd_sc_hd__inv_2
XFILLER_57_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1611_ _1599_/X _1600_/A _1610_/Y VGND VGND VPWR VPWR _1612_/A sky130_fd_sc_hd__o21ai_4
X_1473_ _1820_/A _1473_/B _1473_/C VGND VGND VPWR VPWR _1473_/Y sky130_fd_sc_hd__nor3_4
XFILLER_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1542_ _2194_/Q _1526_/A _1535_/X VGND VGND VPWR VPWR _1542_/X sky130_fd_sc_hd__o21a_4
XFILLER_39_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2025_ _2027_/CLK _2001_/Q VGND VGND VPWR VPWR DATA_TO_HASH[6] sky130_fd_sc_hd__dfxtp_4
XFILLER_50_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1809_ _1804_/C _1809_/B VGND VGND VPWR VPWR _2125_/D sky130_fd_sc_hd__xor2_4
XFILLER_49_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1387_ _1405_/A VGND VGND VPWR VPWR _1387_/X sky130_fd_sc_hd__buf_2
X_1525_ _1525_/A VGND VGND VPWR VPWR _1525_/X sky130_fd_sc_hd__buf_2
X_1456_ _1292_/X _1456_/B VGND VGND VPWR VPWR _1457_/A sky130_fd_sc_hd__nor2_4
XFILLER_42_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2008_ _2013_/CLK _2008_/D VGND VGND VPWR VPWR _1449_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_50_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1241_ _2049_/Q _1180_/B VGND VGND VPWR VPWR _1241_/X sky130_fd_sc_hd__or2_4
X_1310_ _1914_/B VGND VGND VPWR VPWR _1886_/B sky130_fd_sc_hd__buf_2
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1172_ _1172_/A VGND VGND VPWR VPWR _1172_/X sky130_fd_sc_hd__buf_2
XFILLER_9_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1439_ _1737_/D VGND VGND VPWR VPWR _1886_/C sky130_fd_sc_hd__inv_2
X_1508_ _1573_/B _2200_/Q _1507_/X VGND VGND VPWR VPWR _2208_/D sky130_fd_sc_hd__o21a_4
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1790_ _1802_/A _2127_/Q VGND VGND VPWR VPWR _1790_/Y sky130_fd_sc_hd__nand2_4
XFILLER_14_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1224_ _1849_/A _1209_/X _1272_/B VGND VGND VPWR VPWR _1224_/X sky130_fd_sc_hd__a21o_4
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1155_ _1154_/X VGND VGND VPWR VPWR _1230_/B sky130_fd_sc_hd__buf_2
X_1086_ _1086_/A VGND VGND VPWR VPWR _1086_/X sky130_fd_sc_hd__buf_2
X_1988_ _2245_/Q _0996_/A _1987_/X VGND VGND VPWR VPWR _1988_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_m1_clk_local clkbuf_2_3_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_2_3_0_m1_clk_local/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_2_0_addressalyzerBlock.SPI_CLK clkbuf_3_2_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_3_2_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1842_ _1842_/A _1841_/Y VGND VGND VPWR VPWR _2110_/D sky130_fd_sc_hd__xnor2_4
X_1911_ _1042_/Y _1909_/X _1905_/X _1163_/Y _1910_/X VGND VGND VPWR VPWR _2082_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_42_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1773_ _2077_/Q _2101_/Q _1857_/B _1857_/C VGND VGND VPWR VPWR _1856_/B sky130_fd_sc_hd__nand4_4
X_2187_ _2016_/CLK _2187_/D VGND VGND VPWR VPWR _2187_/Q sky130_fd_sc_hd__dfxtp_4
X_1207_ _1207_/A _1207_/B _1207_/C _1207_/D VGND VGND VPWR VPWR _1207_/X sky130_fd_sc_hd__and4_4
XFILLER_33_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1069_ _1062_/Y _1128_/B VGND VGND VPWR VPWR _1069_/Y sky130_fd_sc_hd__nand2_4
X_1138_ _1091_/X _1076_/A _1137_/Y VGND VGND VPWR VPWR _1138_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2041_ _2056_/CLK _2042_/Q VGND VGND VPWR VPWR _2041_/Q sky130_fd_sc_hd__dfxtp_4
X_2110_ _2110_/CLK _2110_/D VGND VGND VPWR VPWR _1842_/A sky130_fd_sc_hd__dfxtp_4
X_1825_ _1825_/A _1827_/A VGND VGND VPWR VPWR _1825_/X sky130_fd_sc_hd__and2_4
X_1756_ _1753_/A _1443_/X _1316_/A VGND VGND VPWR VPWR _1756_/Y sky130_fd_sc_hd__nand3_4
XFILLER_38_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1687_ _1681_/A VGND VGND VPWR VPWR _1689_/A sky130_fd_sc_hd__buf_2
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2239_ _2243_/CLK _1041_/Y VGND VGND VPWR VPWR _1028_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_21_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1610_ _1587_/C _1609_/X _1574_/A _1599_/X _1654_/A VGND VGND VPWR VPWR _1610_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1472_ _1817_/B VGND VGND VPWR VPWR _1820_/A sky130_fd_sc_hd__inv_2
X_1541_ _2194_/Q _1525_/A _1540_/X VGND VGND VPWR VPWR _1541_/X sky130_fd_sc_hd__o21a_4
X_2024_ _2181_/CLK _2024_/D VGND VGND VPWR VPWR DATA_TO_HASH[5] sky130_fd_sc_hd__dfxtp_4
X_1808_ _1807_/Y VGND VGND VPWR VPWR _1808_/Y sky130_fd_sc_hd__inv_2
X_1739_ _1739_/A VGND VGND VPWR VPWR _1739_/X sky130_fd_sc_hd__buf_2
XFILLER_45_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1524_ _1526_/A VGND VGND VPWR VPWR _1525_/A sky130_fd_sc_hd__inv_2
X_1386_ _1382_/X _1385_/Y _1175_/A VGND VGND VPWR VPWR _1386_/X sky130_fd_sc_hd__a21o_4
X_1455_ _2193_/Q _0997_/X _1545_/B _1545_/C VGND VGND VPWR VPWR _1546_/A sky130_fd_sc_hd__nand4_4
XFILLER_35_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2007_ _2013_/CLK _2007_/D VGND VGND VPWR VPWR _2007_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_23_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1240_ _1230_/Y _1231_/Y _1239_/Y VGND VGND VPWR VPWR _1240_/Y sky130_fd_sc_hd__a21oi_4
X_1171_ _1171_/A VGND VGND VPWR VPWR _1171_/X sky130_fd_sc_hd__buf_2
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1507_ _1503_/X _1892_/A _1935_/B VGND VGND VPWR VPWR _1507_/X sky130_fd_sc_hd__o21a_4
XFILLER_55_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1369_ _1369_/A _1397_/B _1369_/C VGND VGND VPWR VPWR _1369_/Y sky130_fd_sc_hd__nand3_4
XFILLER_46_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1438_ _1438_/A _1451_/B _1449_/C VGND VGND VPWR VPWR _1438_/Y sky130_fd_sc_hd__nor3_4
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1154_ _1347_/A VGND VGND VPWR VPWR _1154_/X sky130_fd_sc_hd__buf_2
X_1223_ _1223_/A _1222_/Y VGND VGND VPWR VPWR _1272_/B sky130_fd_sc_hd__nand2_4
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1085_ _1149_/A VGND VGND VPWR VPWR _1104_/A sky130_fd_sc_hd__inv_2
X_1987_ _2246_/Q _1016_/B VGND VGND VPWR VPWR _1987_/X sky130_fd_sc_hd__or2_4
XFILLER_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1910_ _1897_/C _1196_/X _1195_/X _1740_/X _1038_/X VGND VGND VPWR VPWR _1910_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1841_ _2109_/Q _1779_/B _1829_/B _1836_/B VGND VGND VPWR VPWR _1841_/Y sky130_fd_sc_hd__nand4_4
X_1772_ _1772_/A _2103_/Q VGND VGND VPWR VPWR _1774_/C sky130_fd_sc_hd__nand2_4
XFILLER_6_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2186_ _2127_/CLK _1572_/Y VGND VGND VPWR VPWR _2186_/Q sky130_fd_sc_hd__dfxtp_4
X_1206_ _1909_/A VGND VGND VPWR VPWR _1207_/B sky130_fd_sc_hd__inv_2
X_1137_ _1091_/X _1104_/Y _1090_/C _1084_/A _1092_/X VGND VGND VPWR VPWR _1137_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1068_ _1067_/Y VGND VGND VPWR VPWR _1128_/B sky130_fd_sc_hd__inv_2
XFILLER_0_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2040_ _2181_/CLK _1872_/C VGND VGND VPWR VPWR _2034_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_62_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1824_ _2117_/Q _1824_/B VGND VGND VPWR VPWR _1824_/Y sky130_fd_sc_hd__xnor2_4
X_1755_ _1739_/X _1753_/Y _1754_/Y VGND VGND VPWR VPWR _2135_/D sky130_fd_sc_hd__o21ai_4
X_1686_ _1697_/A _2246_/Q VGND VGND VPWR VPWR _2157_/D sky130_fd_sc_hd__and2_4
X_2238_ _2225_/CLK _2238_/D VGND VGND VPWR VPWR _1969_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_38_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2169_ _2173_/CLK _2169_/D VGND VGND VPWR VPWR _1579_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_13_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1540_ _2195_/Q _1526_/A _1535_/X VGND VGND VPWR VPWR _1540_/X sky130_fd_sc_hd__o21a_4
X_1471_ _2127_/Q _1189_/A _1191_/A _1377_/A _1198_/A VGND VGND VPWR VPWR _1471_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2023_ _2127_/CLK _1999_/Q VGND VGND VPWR VPWR DATA_TO_HASH[4] sky130_fd_sc_hd__dfxtp_4
XFILLER_62_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1807_ _1789_/X _1788_/Y VGND VGND VPWR VPWR _1807_/Y sky130_fd_sc_hd__xnor2_4
X_1738_ _1738_/A VGND VGND VPWR VPWR _1739_/A sky130_fd_sc_hd__inv_2
X_1669_ _1581_/B VGND VGND VPWR VPWR _1670_/B sky130_fd_sc_hd__buf_2
XFILLER_26_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1454_ _1454_/A VGND VGND VPWR VPWR _1454_/Y sky130_fd_sc_hd__inv_2
X_1523_ _1501_/Y _2194_/Q _1522_/X VGND VGND VPWR VPWR _1523_/X sky130_fd_sc_hd__o21a_4
X_1385_ _1383_/Y _1233_/X _1384_/Y VGND VGND VPWR VPWR _1385_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_27_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2006_ _2013_/CLK _1961_/Y VGND VGND VPWR VPWR _1309_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_2_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1170_ _1170_/A VGND VGND VPWR VPWR _1170_/X sky130_fd_sc_hd__buf_2
XFILLER_64_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1506_ _1573_/B _2201_/Q _1505_/X VGND VGND VPWR VPWR _1506_/X sky130_fd_sc_hd__o21a_4
X_1437_ _1451_/C VGND VGND VPWR VPWR _1449_/C sky130_fd_sc_hd__inv_2
Xclkbuf_4_2_0_addressalyzerBlock.SPI_CLK clkbuf_4_3_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2202_/CLK sky130_fd_sc_hd__clkbuf_1
X_1368_ _1419_/A _1842_/A _1419_/C VGND VGND VPWR VPWR _1369_/C sky130_fd_sc_hd__nand3_4
X_1299_ _1325_/A _1278_/B _1894_/A VGND VGND VPWR VPWR _1299_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_7_0_addressalyzerBlock.SPI_CLK clkbuf_2_3_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1153_ _1377_/A _1153_/B VGND VGND VPWR VPWR _1153_/Y sky130_fd_sc_hd__nor2_4
X_1222_ _1217_/X _1708_/C _1708_/A VGND VGND VPWR VPWR _1222_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_37_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1084_ _1084_/A VGND VGND VPWR VPWR _1087_/A sky130_fd_sc_hd__inv_2
X_1986_ _2041_/Q _2159_/Q VGND VGND VPWR VPWR IRQ_OUT_toHost sky130_fd_sc_hd__or2_4
XFILLER_20_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1840_ _1838_/A _1838_/B VGND VGND VPWR VPWR _2111_/D sky130_fd_sc_hd__xor2_4
XFILLER_42_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1771_ _1833_/A _2113_/Q VGND VGND VPWR VPWR _1771_/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1205_ _1205_/A _2220_/Q VGND VGND VPWR VPWR _1909_/A sky130_fd_sc_hd__nand2_4
X_2185_ _2202_/CLK _2185_/D VGND VGND VPWR VPWR _1280_/A sky130_fd_sc_hd__dfxtp_4
X_1067_ _1282_/A _1066_/A _1318_/A VGND VGND VPWR VPWR _1067_/Y sky130_fd_sc_hd__nand3_4
X_1136_ _1132_/Y _1134_/Y _1135_/X VGND VGND VPWR VPWR _2232_/D sky130_fd_sc_hd__a21oi_4
X_1969_ _1746_/B _1969_/B _1036_/B _1325_/X VGND VGND VPWR VPWR _1969_/Y sky130_fd_sc_hd__nand4_4
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1823_ _1827_/B _2116_/Q _1827_/A VGND VGND VPWR VPWR _1824_/B sky130_fd_sc_hd__nand3_4
X_1754_ _1763_/A _1757_/B _1460_/A VGND VGND VPWR VPWR _1754_/Y sky130_fd_sc_hd__nand3_4
X_1685_ _1697_/A IRQ_OUT_fromClient VGND VGND VPWR VPWR _1685_/X sky130_fd_sc_hd__and2_4
XFILLER_38_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2237_ _2225_/CLK _1082_/Y VGND VGND VPWR VPWR _1484_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_53_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2099_ _2110_/CLK _2099_/D VGND VGND VPWR VPWR _1857_/C sky130_fd_sc_hd__dfxtp_4
X_2168_ _2173_/CLK _2168_/D VGND VGND VPWR VPWR _1648_/A sky130_fd_sc_hd__dfxtp_4
X_1119_ _1316_/A _1966_/B _1079_/X VGND VGND VPWR VPWR _1119_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_48_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1470_ _1461_/X _1468_/Y _1469_/Y VGND VGND VPWR VPWR _1470_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_39_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2022_ _2022_/CLK _1998_/Q VGND VGND VPWR VPWR DATA_TO_HASH[3] sky130_fd_sc_hd__dfxtp_4
XFILLER_35_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1806_ _1805_/X VGND VGND VPWR VPWR _1806_/Y sky130_fd_sc_hd__inv_2
X_1737_ _1218_/X _1914_/B _1312_/A _1737_/D VGND VGND VPWR VPWR _1738_/A sky130_fd_sc_hd__and4_4
X_1668_ _2162_/Q VGND VGND VPWR VPWR _1678_/B sky130_fd_sc_hd__buf_2
X_1599_ _2181_/Q VGND VGND VPWR VPWR _1599_/X sky130_fd_sc_hd__buf_2
XFILLER_38_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1453_ _1450_/X _1451_/Y _1452_/Y VGND VGND VPWR VPWR _1454_/A sky130_fd_sc_hd__o21ai_4
XFILLER_4_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1522_ _1503_/A _1907_/A _1521_/X VGND VGND VPWR VPWR _1522_/X sky130_fd_sc_hd__o21a_4
XFILLER_55_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1384_ _1164_/X _1879_/C _1172_/X VGND VGND VPWR VPWR _1384_/Y sky130_fd_sc_hd__a21oi_4
X_2005_ _2013_/CLK _2005_/D VGND VGND VPWR VPWR _2005_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_35_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1367_ _1202_/A VGND VGND VPWR VPWR _1419_/C sky130_fd_sc_hd__buf_2
XFILLER_28_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1436_ _1436_/A _1451_/A _1445_/B VGND VGND VPWR VPWR _1436_/Y sky130_fd_sc_hd__nor3_4
X_1505_ _1503_/X _1741_/C _1935_/B VGND VGND VPWR VPWR _1505_/X sky130_fd_sc_hd__o21a_4
X_1298_ _1050_/Y _1104_/A _1298_/C VGND VGND VPWR VPWR _1298_/Y sky130_fd_sc_hd__nand3_4
XFILLER_11_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1221_ _1220_/X VGND VGND VPWR VPWR _1708_/A sky130_fd_sc_hd__buf_2
XFILLER_6_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1152_ _1215_/A _1207_/C _1207_/D _1152_/D VGND VGND VPWR VPWR _1153_/B sky130_fd_sc_hd__nand4_4
XFILLER_37_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1083_ _1147_/B VGND VGND VPWR VPWR _1084_/A sky130_fd_sc_hd__buf_2
X_1985_ _1499_/B MISO_fromClient _1984_/Y VGND VGND VPWR VPWR MISO_toHost sky130_fd_sc_hd__o21a_4
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1419_ _1419_/A _2108_/Q _1419_/C VGND VGND VPWR VPWR _1420_/C sky130_fd_sc_hd__nand3_4
XFILLER_28_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1770_ _1839_/A _1770_/B VGND VGND VPWR VPWR _1831_/A sky130_fd_sc_hd__nand2_4
X_1204_ _1048_/A _1152_/D VGND VGND VPWR VPWR _1207_/A sky130_fd_sc_hd__nor2_4
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2184_ _2022_/CLK _1598_/Y VGND VGND VPWR VPWR CLK_LED sky130_fd_sc_hd__dfxtp_4
X_1066_ _1066_/A _1054_/Y _1066_/C _1066_/D VGND VGND VPWR VPWR _1318_/A sky130_fd_sc_hd__nand4_4
X_1135_ _1070_/X _1482_/B _1446_/A VGND VGND VPWR VPWR _1135_/X sky130_fd_sc_hd__a21o_4
X_1899_ _1898_/Y _1899_/B _1999_/D VGND VGND VPWR VPWR _1899_/Y sky130_fd_sc_hd__nand3_4
X_1968_ _1036_/B _1964_/B _1696_/A _1449_/Y VGND VGND VPWR VPWR _1968_/X sky130_fd_sc_hd__a211o_4
XFILLER_56_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1822_ _1781_/A _1822_/B VGND VGND VPWR VPWR _2118_/D sky130_fd_sc_hd__xor2_4
XFILLER_30_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1753_ _1753_/A _1443_/X _1753_/C VGND VGND VPWR VPWR _1753_/Y sky130_fd_sc_hd__nand3_4
XFILLER_15_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1684_ _1681_/A VGND VGND VPWR VPWR _1697_/A sky130_fd_sc_hd__buf_2
X_2167_ _2173_/CLK _2167_/D VGND VGND VPWR VPWR _1580_/B sky130_fd_sc_hd__dfxtp_4
X_2236_ _2202_/CLK _2236_/D VGND VGND VPWR VPWR _1058_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2098_ _2137_/CLK _1868_/Y VGND VGND VPWR VPWR _2098_/Q sky130_fd_sc_hd__dfxtp_4
X_1049_ _1048_/Y VGND VGND VPWR VPWR _1049_/X sky130_fd_sc_hd__buf_2
XFILLER_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1118_ _1120_/A _1116_/X _1117_/Y VGND VGND VPWR VPWR _1118_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_21_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2021_ _2027_/CLK _1997_/Q VGND VGND VPWR VPWR DATA_TO_HASH[2] sky130_fd_sc_hd__dfxtp_4
XFILLER_50_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1805_ _2127_/Q _1804_/Y VGND VGND VPWR VPWR _1805_/X sky130_fd_sc_hd__xor2_4
X_1736_ _1734_/Y _1213_/A _1735_/Y VGND VGND VPWR VPWR _1736_/Y sky130_fd_sc_hd__a21oi_4
X_1667_ _1661_/A _1661_/B _1666_/Y VGND VGND VPWR VPWR _1667_/Y sky130_fd_sc_hd__a21oi_4
X_1598_ _1597_/Y VGND VGND VPWR VPWR _1598_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2219_ _2050_/CLK _1375_/Y VGND VGND VPWR VPWR _2219_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1383_ _2085_/Q VGND VGND VPWR VPWR _1383_/Y sky130_fd_sc_hd__inv_2
X_1452_ _1450_/X _1480_/A _1293_/X VGND VGND VPWR VPWR _1452_/Y sky130_fd_sc_hd__a21oi_4
X_1521_ _1504_/A VGND VGND VPWR VPWR _1521_/X sky130_fd_sc_hd__buf_2
X_2004_ _2050_/CLK _2003_/Q VGND VGND VPWR VPWR _2004_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_35_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_7_0_addressalyzerBlock.SPI_CLK clkbuf_4_7_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2056_/CLK sky130_fd_sc_hd__clkbuf_1
X_1719_ _2059_/Q VGND VGND VPWR VPWR _1720_/B sky130_fd_sc_hd__inv_2
XFILLER_58_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1504_ _1504_/A VGND VGND VPWR VPWR _1935_/B sky130_fd_sc_hd__buf_2
X_1366_ _1366_/A VGND VGND VPWR VPWR _1419_/A sky130_fd_sc_hd__inv_2
X_1435_ _1438_/A VGND VGND VPWR VPWR _1445_/B sky130_fd_sc_hd__inv_2
X_1297_ _1296_/Y _1282_/A _1318_/A _1282_/C _1104_/A VGND VGND VPWR VPWR _1297_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_46_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1220_ _1207_/A _1207_/C _1207_/D VGND VGND VPWR VPWR _1220_/X sky130_fd_sc_hd__and3_4
X_1151_ _1184_/A VGND VGND VPWR VPWR _1152_/D sky130_fd_sc_hd__inv_2
X_1082_ _1077_/Y _1080_/Y _1081_/Y VGND VGND VPWR VPWR _1082_/Y sky130_fd_sc_hd__a21oi_4
X_1984_ _1983_/Y _1499_/B VGND VGND VPWR VPWR _1984_/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1418_ _1403_/Y _1416_/Y _1417_/X VGND VGND VPWR VPWR _1420_/A sky130_fd_sc_hd__o21ai_4
X_1349_ _1405_/A _1348_/Y VGND VGND VPWR VPWR _1349_/Y sky130_fd_sc_hd__nor2_4
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1203_ _1202_/Y _1198_/A VGND VGND VPWR VPWR _1203_/Y sky130_fd_sc_hd__nor2_4
X_2183_ _2022_/CLK _1603_/X VGND VGND VPWR VPWR _1596_/C sky130_fd_sc_hd__dfxtp_4
X_1134_ _1762_/C _1123_/X _1079_/X VGND VGND VPWR VPWR _1134_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_33_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1065_ _2005_/Q VGND VGND VPWR VPWR _1066_/C sky130_fd_sc_hd__inv_2
XFILLER_18_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1898_ _1897_/X VGND VGND VPWR VPWR _1898_/Y sky130_fd_sc_hd__inv_2
X_1967_ _1282_/C _1966_/Y _1446_/X VGND VGND VPWR VPWR _2009_/D sky130_fd_sc_hd__a21oi_4
XFILLER_0_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1821_ _1825_/A _2117_/Q _2116_/Q _1827_/A VGND VGND VPWR VPWR _1822_/B sky130_fd_sc_hd__and4_4
X_1752_ _1739_/X _1932_/A _1751_/Y VGND VGND VPWR VPWR _1752_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_30_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1683_ _1701_/A _2158_/Q VGND VGND VPWR VPWR _2159_/D sky130_fd_sc_hd__and2_4
XFILLER_57_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2097_ _2137_/CLK _2097_/D VGND VGND VPWR VPWR _2097_/Q sky130_fd_sc_hd__dfxtp_4
X_2166_ _2173_/CLK _1667_/Y VGND VGND VPWR VPWR _1660_/A sky130_fd_sc_hd__dfxtp_4
X_2235_ _2225_/CLK _2235_/D VGND VGND VPWR VPWR _1057_/A sky130_fd_sc_hd__dfxtp_4
X_1117_ _1120_/A _1106_/X _1126_/A _1116_/C _1092_/X VGND VGND VPWR VPWR _1117_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1048_ _1048_/A _1914_/B _1311_/A _2220_/Q VGND VGND VPWR VPWR _1048_/Y sky130_fd_sc_hd__nand4_4
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2020_ _2016_/CLK _1996_/Q VGND VGND VPWR VPWR DATA_TO_HASH[1] sky130_fd_sc_hd__dfxtp_4
XFILLER_62_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1804_ _1804_/A _1804_/B _1804_/C _2124_/Q VGND VGND VPWR VPWR _1804_/Y sky130_fd_sc_hd__nand4_4
X_1735_ _1213_/A _2139_/Q VGND VGND VPWR VPWR _1735_/Y sky130_fd_sc_hd__nor2_4
X_1666_ _1661_/A _1661_/B _1746_/B VGND VGND VPWR VPWR _1666_/Y sky130_fd_sc_hd__o21ai_4
X_1597_ _1591_/Y _1307_/B _1596_/Y VGND VGND VPWR VPWR _1597_/Y sky130_fd_sc_hd__nand3_4
X_2218_ _2243_/CLK _2218_/D VGND VGND VPWR VPWR _1400_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_26_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2149_ _2153_/CLK _1698_/X VGND VGND VPWR VPWR _2149_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_5_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0_m1_clk_local clkbuf_0_m1_clk_local/X VGND VGND VPWR VPWR clkbuf_2_3_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1520_ _1501_/Y _2195_/Q _1519_/X VGND VGND VPWR VPWR _1520_/X sky130_fd_sc_hd__o21a_4
X_1382_ _1922_/C _1154_/X _1166_/X _1381_/Y VGND VGND VPWR VPWR _1382_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_4_12_0_addressalyzerBlock.SPI_CLK clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2214_/CLK sky130_fd_sc_hd__clkbuf_1
X_1451_ _1451_/A _1451_/B _1451_/C VGND VGND VPWR VPWR _1451_/Y sky130_fd_sc_hd__nor3_4
XFILLER_50_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2003_ _2050_/CLK _2003_/D VGND VGND VPWR VPWR _2003_/Q sky130_fd_sc_hd__dfxtp_4
X_1718_ _1718_/A _1718_/B VGND VGND VPWR VPWR _1718_/Y sky130_fd_sc_hd__nand2_4
X_1649_ _1647_/Y _1648_/X _1643_/X _1644_/X VGND VGND VPWR VPWR _1649_/X sky130_fd_sc_hd__and4_4
XFILLER_58_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1503_ _1503_/A VGND VGND VPWR VPWR _1503_/X sky130_fd_sc_hd__buf_2
XFILLER_55_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1365_ _1365_/A VGND VGND VPWR VPWR _1397_/B sky130_fd_sc_hd__buf_2
X_1434_ _1426_/Y _1430_/Y _1433_/X VGND VGND VPWR VPWR _2216_/D sky130_fd_sc_hd__a21oi_4
X_1296_ _1086_/X _1049_/X _1056_/Y VGND VGND VPWR VPWR _1296_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_31_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1150_ _1150_/A VGND VGND VPWR VPWR _1207_/D sky130_fd_sc_hd__buf_2
Xclkbuf_3_4_0_m1_clk_local clkbuf_3_4_0_m1_clk_local/A VGND VGND VPWR VPWR _2110_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1081_ _1484_/A _1128_/B _1031_/X VGND VGND VPWR VPWR _1081_/Y sky130_fd_sc_hd__o21ai_4
X_1983_ _2157_/Q VGND VGND VPWR VPWR _1983_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1417_ _1313_/C _2116_/Q _1313_/B _1366_/A VGND VGND VPWR VPWR _1417_/X sky130_fd_sc_hd__a211o_4
X_1348_ _2070_/Q VGND VGND VPWR VPWR _1348_/Y sky130_fd_sc_hd__inv_2
X_1279_ _1279_/A VGND VGND VPWR VPWR _1279_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1202_ _1202_/A VGND VGND VPWR VPWR _1202_/Y sky130_fd_sc_hd__inv_2
X_1064_ _1325_/A VGND VGND VPWR VPWR _1066_/A sky130_fd_sc_hd__inv_2
X_2182_ _2181_/CLK _1606_/X VGND VGND VPWR VPWR _1589_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1133_ _1904_/A VGND VGND VPWR VPWR _1762_/C sky130_fd_sc_hd__buf_2
X_1966_ _1036_/B _1966_/B VGND VGND VPWR VPWR _1966_/Y sky130_fd_sc_hd__nand2_4
XFILLER_18_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1897_ _1217_/X _1934_/A _1897_/C VGND VGND VPWR VPWR _1897_/X sky130_fd_sc_hd__and3_4
XFILLER_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1820_ _1820_/A _1820_/B VGND VGND VPWR VPWR _2119_/D sky130_fd_sc_hd__xor2_4
X_1751_ _1763_/A _1757_/B _1253_/A VGND VGND VPWR VPWR _1751_/Y sky130_fd_sc_hd__nand3_4
X_1682_ _1701_/A _1682_/B VGND VGND VPWR VPWR _1682_/X sky130_fd_sc_hd__and2_4
X_2234_ _2202_/CLK _2234_/D VGND VGND VPWR VPWR _1057_/B sky130_fd_sc_hd__dfxtp_4
X_1047_ _1205_/A VGND VGND VPWR VPWR _1311_/A sky130_fd_sc_hd__buf_2
X_2096_ _2207_/CLK _2096_/D VGND VGND VPWR VPWR _1872_/C sky130_fd_sc_hd__dfxtp_4
X_2165_ _2173_/CLK _1673_/X VGND VGND VPWR VPWR _1581_/D sky130_fd_sc_hd__dfxtp_4
X_1116_ _1052_/X _1126_/A _1116_/C _1090_/B VGND VGND VPWR VPWR _1116_/X sky130_fd_sc_hd__and4_4
X_1949_ _1948_/X VGND VGND VPWR VPWR _1949_/X sky130_fd_sc_hd__buf_2
XFILLER_21_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1803_ _1803_/A _1787_/Y VGND VGND VPWR VPWR _1804_/B sky130_fd_sc_hd__nor2_4
XFILLER_50_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1734_ _1709_/X _1731_/Y _1733_/X VGND VGND VPWR VPWR _1734_/Y sky130_fd_sc_hd__o21ai_4
X_1665_ _1917_/A VGND VGND VPWR VPWR _1746_/B sky130_fd_sc_hd__buf_2
X_1596_ _1596_/A _1596_/B _1596_/C CLK_LED VGND VGND VPWR VPWR _1596_/Y sky130_fd_sc_hd__nand4_4
XFILLER_58_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2217_ _2050_/CLK _2217_/D VGND VGND VPWR VPWR _1424_/B sky130_fd_sc_hd__dfxtp_4
X_2079_ _2069_/CLK _1919_/Y VGND VGND VPWR VPWR _1918_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_41_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2148_ _2216_/CLK _2148_/D VGND VGND VPWR VPWR _2148_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_30_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1450_ _1438_/A _1092_/A _1448_/Y _1449_/Y VGND VGND VPWR VPWR _1450_/X sky130_fd_sc_hd__a211o_4
X_1381_ _1405_/A _1380_/Y VGND VGND VPWR VPWR _1381_/Y sky130_fd_sc_hd__nor2_4
XFILLER_50_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2002_ _2022_/CLK _2090_/Q VGND VGND VPWR VPWR _2026_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_23_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1717_ _1715_/Y _1170_/X _1716_/Y VGND VGND VPWR VPWR _1718_/B sky130_fd_sc_hd__o21ai_4
X_1648_ _1648_/A VGND VGND VPWR VPWR _1648_/X sky130_fd_sc_hd__buf_2
X_1579_ _1579_/A VGND VGND VPWR VPWR _1582_/B sky130_fd_sc_hd__inv_2
XFILLER_58_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1433_ _1429_/X _1432_/Y _1293_/X VGND VGND VPWR VPWR _1433_/X sky130_fd_sc_hd__a21o_4
X_1502_ _1501_/Y VGND VGND VPWR VPWR _1573_/B sky130_fd_sc_hd__buf_2
XFILLER_48_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1364_ _1346_/X _1361_/Y _1363_/X VGND VGND VPWR VPWR _1369_/A sky130_fd_sc_hd__o21ai_4
X_1295_ _1289_/Y _1290_/Y _1294_/X VGND VGND VPWR VPWR _1295_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_46_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_3_0_addressalyzerBlock.SPI_CLK clkbuf_2_3_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_2_3_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1080_ _1892_/A _1966_/B _1079_/X VGND VGND VPWR VPWR _1080_/Y sky130_fd_sc_hd__a21oi_4
X_1982_ _1980_/Y S1_CLK_SELECT _1981_/Y VGND VGND VPWR VPWR _1982_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_9_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1416_ _1414_/Y _1285_/X _1415_/Y VGND VGND VPWR VPWR _1416_/Y sky130_fd_sc_hd__a21oi_4
X_1347_ _1347_/A VGND VGND VPWR VPWR _1405_/A sky130_fd_sc_hd__buf_2
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1278_ _1325_/A _1278_/B VGND VGND VPWR VPWR _1279_/A sky130_fd_sc_hd__nor2_4
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1201_ _1311_/A _1312_/A VGND VGND VPWR VPWR _1202_/A sky130_fd_sc_hd__nor2_4
X_2181_ _2181_/CLK _1612_/Y VGND VGND VPWR VPWR _2181_/Q sky130_fd_sc_hd__dfxtp_4
X_1063_ _1092_/A _1066_/D _1280_/A VGND VGND VPWR VPWR _1282_/A sky130_fd_sc_hd__a21o_4
X_1132_ _1116_/C _1106_/X _1129_/Y VGND VGND VPWR VPWR _1132_/Y sky130_fd_sc_hd__o21ai_4
X_1965_ _1964_/Y _1445_/C _1446_/X VGND VGND VPWR VPWR _1965_/Y sky130_fd_sc_hd__a21oi_4
X_1896_ _1886_/A _1886_/C VGND VGND VPWR VPWR _1934_/A sky130_fd_sc_hd__nor2_4
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1750_ _1750_/A VGND VGND VPWR VPWR _1757_/B sky130_fd_sc_hd__buf_2
X_1681_ _1681_/A VGND VGND VPWR VPWR _1701_/A sky130_fd_sc_hd__buf_2
XFILLER_38_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2164_ _2173_/CLK _2164_/D VGND VGND VPWR VPWR _2164_/Q sky130_fd_sc_hd__dfxtp_4
X_2233_ _2225_/CLK _1131_/Y VGND VGND VPWR VPWR _1057_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_53_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1046_ _1184_/A VGND VGND VPWR VPWR _1914_/B sky130_fd_sc_hd__buf_2
X_2095_ _2137_/CLK _2095_/D VGND VGND VPWR VPWR _2039_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1115_ _1963_/A _1115_/B VGND VGND VPWR VPWR _2235_/D sky130_fd_sc_hd__nor2_4
X_1948_ _1218_/X _1144_/B _1886_/B _1927_/D _1292_/X VGND VGND VPWR VPWR _1948_/X
+ sky130_fd_sc_hd__a41o_4
X_1879_ _1874_/A _1899_/B _1879_/C VGND VGND VPWR VPWR _1879_/Y sky130_fd_sc_hd__nand3_4
XFILLER_21_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1802_ _1802_/A _1801_/Y VGND VGND VPWR VPWR _2128_/D sky130_fd_sc_hd__xnor2_4
X_1733_ _1215_/A _2041_/Q _1215_/B _1732_/X VGND VGND VPWR VPWR _1733_/X sky130_fd_sc_hd__or4_4
X_1664_ _1663_/X VGND VGND VPWR VPWR _2167_/D sky130_fd_sc_hd__inv_2
X_1595_ _1574_/Y _1595_/B _1595_/C VGND VGND VPWR VPWR _1596_/B sky130_fd_sc_hd__nor3_4
X_2147_ _2216_/CLK _2147_/D VGND VGND VPWR VPWR _2147_/Q sky130_fd_sc_hd__dfxtp_4
X_2216_ _2216_/CLK _2216_/D VGND VGND VPWR VPWR _2216_/Q sky130_fd_sc_hd__dfxtp_4
X_2078_ _2069_/CLK _1921_/Y VGND VGND VPWR VPWR HASH_LED sky130_fd_sc_hd__dfxtp_4
XFILLER_14_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1029_ _2240_/Q _0997_/X _1028_/X VGND VGND VPWR VPWR _1029_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_39_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1380_ _1380_/A VGND VGND VPWR VPWR _1380_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2001_ _2027_/CLK _2089_/Q VGND VGND VPWR VPWR _2001_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1716_ _1170_/A _1883_/C _1172_/A VGND VGND VPWR VPWR _1716_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_58_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1578_ _1648_/A VGND VGND VPWR VPWR _1582_/A sky130_fd_sc_hd__inv_2
X_1647_ _1647_/A _1661_/B VGND VGND VPWR VPWR _1647_/Y sky130_fd_sc_hd__nor2_4
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1363_ _1313_/C _1781_/A _1313_/B _1366_/A VGND VGND VPWR VPWR _1363_/X sky130_fd_sc_hd__a211o_4
X_1432_ _1971_/A _1971_/C _1066_/C VGND VGND VPWR VPWR _1432_/Y sky130_fd_sc_hd__nand3_4
X_1501_ _1503_/A VGND VGND VPWR VPWR _1501_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1294_ _1339_/A _1087_/A _1293_/X VGND VGND VPWR VPWR _1294_/X sky130_fd_sc_hd__a21o_4
XFILLER_54_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1981_ _1981_/A S1_CLK_SELECT VGND VGND VPWR VPWR _1981_/Y sky130_fd_sc_hd__nor2_4
XFILLER_9_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1415_ _1180_/B _2044_/Q _1188_/A VGND VGND VPWR VPWR _1415_/Y sky130_fd_sc_hd__o21ai_4
X_1346_ _1187_/A _1804_/A _1153_/Y VGND VGND VPWR VPWR _1346_/X sky130_fd_sc_hd__a21o_4
XFILLER_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1277_ _1090_/C _1087_/Y _1276_/Y VGND VGND VPWR VPWR _1277_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_51_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1200_ _1153_/Y _1193_/Y _1199_/X VGND VGND VPWR VPWR _1200_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_2_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2180_ _2181_/CLK _1614_/Y VGND VGND VPWR VPWR _1574_/A sky130_fd_sc_hd__dfxtp_4
X_1131_ _1128_/Y _1130_/Y _1040_/X VGND VGND VPWR VPWR _1131_/Y sky130_fd_sc_hd__a21oi_4
X_1062_ _1042_/Y _1066_/D _1061_/Y VGND VGND VPWR VPWR _1062_/Y sky130_fd_sc_hd__o21ai_4
X_1895_ _1894_/Y _1885_/X _1888_/X _1258_/Y _1890_/X VGND VGND VPWR VPWR _2088_/D
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_3_0_0_m1_clk_local clkbuf_3_1_0_m1_clk_local/A VGND VGND VPWR VPWR _2181_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_1964_ _1964_/A _1964_/B VGND VGND VPWR VPWR _1964_/Y sky130_fd_sc_hd__nand2_4
XFILLER_56_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1329_ _1152_/D VGND VGND VPWR VPWR _1897_/C sky130_fd_sc_hd__buf_2
XFILLER_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1680_ _1963_/A _1693_/B VGND VGND VPWR VPWR _1680_/Y sky130_fd_sc_hd__nor2_4
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2163_ _2173_/CLK _2163_/D VGND VGND VPWR VPWR _1581_/B sky130_fd_sc_hd__dfxtp_4
X_1114_ _1057_/A _1111_/X _1113_/Y _1128_/B VGND VGND VPWR VPWR _1115_/B sky130_fd_sc_hd__a22oi_4
X_2232_ _2202_/CLK _2232_/D VGND VGND VPWR VPWR _1124_/A sky130_fd_sc_hd__dfxtp_4
X_1045_ _1149_/B VGND VGND VPWR VPWR _1086_/A sky130_fd_sc_hd__inv_2
X_2094_ _2137_/CLK _2094_/D VGND VGND VPWR VPWR _2094_/Q sky130_fd_sc_hd__dfxtp_4
X_1947_ _1892_/Y _1944_/A _1946_/Y VGND VGND VPWR VPWR _1947_/Y sky130_fd_sc_hd__o21ai_4
X_1878_ _1756_/Y _1865_/X _1877_/Y VGND VGND VPWR VPWR _2094_/D sky130_fd_sc_hd__o21ai_4
XFILLER_56_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1801_ _2127_/Q _1809_/B _1789_/X _1804_/C VGND VGND VPWR VPWR _1801_/Y sky130_fd_sc_hd__nand4_4
X_1732_ _1732_/A VGND VGND VPWR VPWR _1732_/X sky130_fd_sc_hd__buf_2
X_1663_ _1580_/B _1661_/Y _1662_/Y VGND VGND VPWR VPWR _1663_/X sky130_fd_sc_hd__a21o_4
XFILLER_7_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1594_ _1588_/B VGND VGND VPWR VPWR _1595_/C sky130_fd_sc_hd__buf_2
X_2077_ _2077_/CLK _1923_/Y VGND VGND VPWR VPWR _2077_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2215_ _2077_/CLK _1447_/Y VGND VGND VPWR VPWR _1737_/D sky130_fd_sc_hd__dfxtp_4
X_2146_ _2153_/CLK _1701_/Y VGND VGND VPWR VPWR _2146_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1028_ _1028_/A _0996_/A VGND VGND VPWR VPWR _1028_/X sky130_fd_sc_hd__or2_4
XFILLER_30_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2000_ _2181_/CLK _1258_/A VGND VGND VPWR VPWR _2024_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_3_3_0_addressalyzerBlock.SPI_CLK clkbuf_3_2_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR clkbuf_4_7_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_50_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1715_ _1715_/A VGND VGND VPWR VPWR _1715_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1646_ _1645_/X _1307_/B _1646_/C VGND VGND VPWR VPWR _1646_/X sky130_fd_sc_hd__and3_4
XFILLER_58_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1577_ _1577_/A VGND VGND VPWR VPWR _1577_/Y sky130_fd_sc_hd__inv_2
X_2129_ _2127_/CLK _2129_/D VGND VGND VPWR VPWR _2129_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1500_ _1498_/Y _1499_/Y _1446_/X VGND VGND VPWR VPWR _2210_/D sky130_fd_sc_hd__a21oi_4
XFILLER_9_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1362_ _1198_/A VGND VGND VPWR VPWR _1366_/A sky130_fd_sc_hd__buf_2
X_1431_ _2007_/Q VGND VGND VPWR VPWR _1971_/C sky130_fd_sc_hd__inv_2
X_1293_ _1292_/X VGND VGND VPWR VPWR _1293_/X sky130_fd_sc_hd__buf_2
XFILLER_51_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1629_ _1628_/Y VGND VGND VPWR VPWR _2177_/D sky130_fd_sc_hd__inv_2
XFILLER_39_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1980_ S1_CLK_IN VGND VGND VPWR VPWR _1980_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1414_ _1414_/A _1413_/X VGND VGND VPWR VPWR _1414_/Y sky130_fd_sc_hd__nand2_4
X_1345_ _1344_/X VGND VGND VPWR VPWR _1345_/X sky130_fd_sc_hd__buf_2
XFILLER_28_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1276_ _1090_/C _1050_/Y _1084_/A _1149_/A _1092_/X VGND VGND VPWR VPWR _1276_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_51_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1130_ _1070_/X _1129_/Y _1126_/A VGND VGND VPWR VPWR _1130_/Y sky130_fd_sc_hd__o21ai_4
X_1061_ _1061_/A _1076_/A _1056_/Y _1061_/D VGND VGND VPWR VPWR _1061_/Y sky130_fd_sc_hd__nand4_4
XFILLER_18_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1894_ _1894_/A VGND VGND VPWR VPWR _1894_/Y sky130_fd_sc_hd__inv_2
X_1963_ _1963_/A _1963_/B VGND VGND VPWR VPWR _2010_/D sky130_fd_sc_hd__nor2_4
X_1259_ _1171_/X _1872_/C _1172_/A VGND VGND VPWR VPWR _1259_/Y sky130_fd_sc_hd__a21oi_4
X_1328_ _1886_/B _1207_/B _1314_/X VGND VGND VPWR VPWR _1328_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2231_ _2225_/CLK _1142_/Y VGND VGND VPWR VPWR _1105_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_53_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2093_ _2137_/CLK _2093_/D VGND VGND VPWR VPWR _1879_/C sky130_fd_sc_hd__dfxtp_4
X_2162_ _2173_/CLK _2162_/D VGND VGND VPWR VPWR _2162_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1044_ _1969_/B VGND VGND VPWR VPWR _1061_/A sky130_fd_sc_hd__inv_2
X_1113_ _1057_/A _1126_/C _1109_/Y _1112_/Y _1066_/D VGND VGND VPWR VPWR _1113_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1946_ _1944_/A _1341_/C _2065_/Q VGND VGND VPWR VPWR _1946_/Y sky130_fd_sc_hd__nand3_4
X_1877_ _1874_/A _1899_/B _2094_/Q VGND VGND VPWR VPWR _1877_/Y sky130_fd_sc_hd__nand3_4
XFILLER_60_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1800_ _1799_/Y VGND VGND VPWR VPWR _2129_/D sky130_fd_sc_hd__inv_2
XFILLER_35_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1731_ _1731_/A _1731_/B VGND VGND VPWR VPWR _1731_/Y sky130_fd_sc_hd__nor2_4
X_1662_ _1580_/B _1661_/Y _1681_/A VGND VGND VPWR VPWR _1662_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_7_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2214_ _2214_/CLK _1454_/Y VGND VGND VPWR VPWR _1213_/A sky130_fd_sc_hd__dfxtp_4
X_1593_ _2181_/Q VGND VGND VPWR VPWR _1595_/B sky130_fd_sc_hd__inv_2
XFILLER_53_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2076_ _2069_/CLK _2076_/D VGND VGND VPWR VPWR _2076_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_41_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2145_ _2153_/CLK _1702_/Y VGND VGND VPWR VPWR _2145_/Q sky130_fd_sc_hd__dfxtp_4
X_1027_ _1025_/Y _1003_/X _1026_/Y VGND VGND VPWR VPWR _1027_/Y sky130_fd_sc_hd__a21oi_4
X_1929_ _1935_/A _1341_/C _2074_/Q _1185_/A _1928_/Y VGND VGND VPWR VPWR _2074_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_55_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1714_ _1712_/Y _1170_/X _1713_/Y VGND VGND VPWR VPWR _1718_/A sky130_fd_sc_hd__o21ai_4
X_1645_ _1642_/Y _1643_/X _1644_/X _1583_/C _2172_/Q VGND VGND VPWR VPWR _1645_/X
+ sky130_fd_sc_hd__a41o_4
X_1576_ _1576_/A VGND VGND VPWR VPWR _1608_/B sky130_fd_sc_hd__inv_2
XFILLER_54_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2128_ _2127_/CLK _2128_/D VGND VGND VPWR VPWR _1802_/A sky130_fd_sc_hd__dfxtp_4
X_2059_ _2142_/CLK _2059_/D VGND VGND VPWR VPWR _2059_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1430_ _1436_/A _1325_/X _2007_/Q _2005_/Q _1429_/X VGND VGND VPWR VPWR _1430_/Y
+ sky130_fd_sc_hd__o41ai_4
X_1361_ _1359_/Y _1285_/X _1360_/Y VGND VGND VPWR VPWR _1361_/Y sky130_fd_sc_hd__a21oi_4
X_1292_ _1886_/A VGND VGND VPWR VPWR _1292_/X sky130_fd_sc_hd__buf_2
XFILLER_23_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1559_ _1981_/A _1565_/A SPI_CLK_RESET_N VGND VGND VPWR VPWR _1559_/Y sky130_fd_sc_hd__o21ai_4
X_1628_ _1628_/A _1628_/B VGND VGND VPWR VPWR _1628_/Y sky130_fd_sc_hd__nand2_4
XFILLER_46_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1413_ _1763_/C _1355_/X _1161_/A _1412_/Y VGND VGND VPWR VPWR _1413_/X sky130_fd_sc_hd__a211o_4
X_1344_ _1708_/C _1207_/A _1207_/C _1207_/D VGND VGND VPWR VPWR _1344_/X sky130_fd_sc_hd__and4_4
X_1275_ _1275_/A _1274_/Y VGND VGND VPWR VPWR _2228_/D sky130_fd_sc_hd__nand2_4
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1060_ _1060_/A VGND VGND VPWR VPWR _1061_/D sky130_fd_sc_hd__buf_2
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1962_ _1456_/B _2005_/Q _1964_/A _1966_/B VGND VGND VPWR VPWR _1963_/B sky130_fd_sc_hd__a22oi_4
X_1893_ _1892_/Y _1885_/X _1888_/X _1236_/Y _1890_/X VGND VGND VPWR VPWR _1893_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_56_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1258_ _1258_/A VGND VGND VPWR VPWR _1258_/Y sky130_fd_sc_hd__inv_2
X_1189_ _1189_/A VGND VGND VPWR VPWR _1265_/B sky130_fd_sc_hd__buf_2
X_1327_ _1325_/X _1123_/X _1902_/A VGND VGND VPWR VPWR _1327_/Y sky130_fd_sc_hd__o21ai_4
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2230_ _2243_/CLK _1229_/Y VGND VGND VPWR VPWR _2230_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2092_ _2137_/CLK _2092_/D VGND VGND VPWR VPWR _2036_/D sky130_fd_sc_hd__dfxtp_4
X_1112_ _1753_/C VGND VGND VPWR VPWR _1112_/Y sky130_fd_sc_hd__inv_2
X_2161_ _2153_/CLK _1680_/Y VGND VGND VPWR VPWR _1693_/D sky130_fd_sc_hd__dfxtp_4
X_1043_ _1278_/B VGND VGND VPWR VPWR _1066_/D sky130_fd_sc_hd__inv_2
X_1945_ _1042_/Y _1944_/A _1944_/Y VGND VGND VPWR VPWR _1945_/Y sky130_fd_sc_hd__o21ai_4
X_1876_ _1750_/A VGND VGND VPWR VPWR _1899_/B sky130_fd_sc_hd__buf_2
XFILLER_56_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_3_0_addressalyzerBlock.SPI_CLK clkbuf_4_3_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2142_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_47_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1730_ _1725_/Y _1727_/X _1729_/Y VGND VGND VPWR VPWR _1731_/B sky130_fd_sc_hd__a21oi_4
X_1661_ _1661_/A _1661_/B VGND VGND VPWR VPWR _1661_/Y sky130_fd_sc_hd__nor2_4
XFILLER_7_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1592_ _1589_/C VGND VGND VPWR VPWR _1596_/A sky130_fd_sc_hd__buf_2
XFILLER_38_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2144_ _2225_/CLK _1703_/X VGND VGND VPWR VPWR _2144_/Q sky130_fd_sc_hd__dfxtp_4
X_2213_ _2202_/CLK _2213_/D VGND VGND VPWR VPWR _1503_/A sky130_fd_sc_hd__dfxtp_4
X_2075_ _2042_/CLK _1926_/Y VGND VGND VPWR VPWR _2015_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_53_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1026_ _1400_/B _1003_/A _1008_/X VGND VGND VPWR VPWR _1026_/Y sky130_fd_sc_hd__o21ai_4
X_1928_ _1928_/A VGND VGND VPWR VPWR _1928_/Y sky130_fd_sc_hd__inv_2
X_1859_ _1858_/X VGND VGND VPWR VPWR _1859_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_2_2_0_m1_clk_local clkbuf_2_3_0_m1_clk_local/A VGND VGND VPWR VPWR clkbuf_3_4_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1713_ _1171_/X _2067_/Q _1166_/A VGND VGND VPWR VPWR _1713_/Y sky130_fd_sc_hd__a21oi_4
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1644_ _1644_/A VGND VGND VPWR VPWR _1644_/X sky130_fd_sc_hd__buf_2
X_1575_ _2173_/Q VGND VGND VPWR VPWR _1575_/Y sky130_fd_sc_hd__inv_2
X_2127_ _2127_/CLK _1806_/Y VGND VGND VPWR VPWR _2127_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_58_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2058_ _2050_/CLK DATA_FROM_HASH[7] VGND VGND VPWR VPWR _2050_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_34_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1009_ _1251_/B _1004_/X _1008_/X VGND VGND VPWR VPWR _1009_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_26_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1360_ _1285_/X _2046_/Q _1188_/X VGND VGND VPWR VPWR _1360_/Y sky130_fd_sc_hd__o21ai_4
X_1291_ _1283_/A VGND VGND VPWR VPWR _1339_/A sky130_fd_sc_hd__buf_2
XFILLER_63_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1558_ _1563_/A _1562_/C _1570_/C VGND VGND VPWR VPWR _1565_/A sky130_fd_sc_hd__nor3_4
X_1489_ _1487_/Y _1057_/A _1120_/A _1357_/B VGND VGND VPWR VPWR _1489_/Y sky130_fd_sc_hd__a22oi_4
X_1627_ _1621_/C _1609_/A _1585_/A _1585_/B VGND VGND VPWR VPWR _1628_/B sky130_fd_sc_hd__nand4_4
XFILLER_54_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1412_ _1387_/X _1412_/B VGND VGND VPWR VPWR _1412_/Y sky130_fd_sc_hd__nor2_4
X_1343_ _1217_/X _1708_/A _1480_/A _1215_/Y VGND VGND VPWR VPWR _1343_/X sky130_fd_sc_hd__a211o_4
XFILLER_51_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1274_ _1274_/A _1274_/B VGND VGND VPWR VPWR _1274_/Y sky130_fd_sc_hd__nand2_4
XFILLER_59_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1892_ _1892_/A VGND VGND VPWR VPWR _1892_/Y sky130_fd_sc_hd__inv_2
X_1961_ _1957_/A _1964_/A _1971_/C _1320_/Y _1960_/X VGND VGND VPWR VPWR _1961_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1326_ _2204_/Q VGND VGND VPWR VPWR _1902_/A sky130_fd_sc_hd__buf_2
X_1188_ _1188_/A VGND VGND VPWR VPWR _1188_/X sky130_fd_sc_hd__buf_2
X_1257_ _1255_/Y _1233_/X _1256_/Y VGND VGND VPWR VPWR _1257_/Y sky130_fd_sc_hd__o21ai_4
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XINSDIODE2_0 ID_fromClient VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2160_ _2153_/CLK _1682_/X VGND VGND VPWR VPWR _2160_/Q sky130_fd_sc_hd__dfxtp_4
X_2091_ _2137_/CLK _1884_/Y VGND VGND VPWR VPWR _1883_/C sky130_fd_sc_hd__dfxtp_4
X_1042_ _1741_/C VGND VGND VPWR VPWR _1042_/Y sky130_fd_sc_hd__inv_2
X_1111_ _1109_/Y _1298_/C _1067_/Y VGND VGND VPWR VPWR _1111_/X sky130_fd_sc_hd__a21o_4
X_1944_ _1944_/A _1918_/B _2066_/Q VGND VGND VPWR VPWR _1944_/Y sky130_fd_sc_hd__nand3_4
X_1875_ _1753_/Y _1865_/X _1874_/Y VGND VGND VPWR VPWR _2095_/D sky130_fd_sc_hd__o21ai_4
XFILLER_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1309_ _1309_/A VGND VGND VPWR VPWR _1451_/A sky130_fd_sc_hd__buf_2
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1660_ _1660_/A VGND VGND VPWR VPWR _1661_/A sky130_fd_sc_hd__inv_2
X_1591_ _1589_/Y _1590_/Y VGND VGND VPWR VPWR _1591_/Y sky130_fd_sc_hd__nand2_4
X_2212_ _2050_/CLK _2212_/D VGND VGND VPWR VPWR _1480_/B sky130_fd_sc_hd__dfxtp_4
X_2143_ _2216_/CLK _2143_/D VGND VGND VPWR VPWR _2143_/Q sky130_fd_sc_hd__dfxtp_4
X_2074_ _2137_/CLK _2074_/D VGND VGND VPWR VPWR _2074_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1025_ _2240_/Q _0996_/A _1024_/X VGND VGND VPWR VPWR _1025_/Y sky130_fd_sc_hd__o21ai_4
X_1858_ _2101_/Q _1857_/Y VGND VGND VPWR VPWR _1858_/X sky130_fd_sc_hd__xor2_4
X_1927_ _1897_/C _1144_/B _1196_/X _1927_/D VGND VGND VPWR VPWR _1935_/A sky130_fd_sc_hd__nand4_4
X_1789_ _1804_/A VGND VGND VPWR VPWR _1789_/X sky130_fd_sc_hd__buf_2
XFILLER_39_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1712_ _2015_/D VGND VGND VPWR VPWR _1712_/Y sky130_fd_sc_hd__inv_2
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1643_ _1579_/A VGND VGND VPWR VPWR _1643_/X sky130_fd_sc_hd__buf_2
XFILLER_6_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1574_ _1574_/A VGND VGND VPWR VPWR _1574_/Y sky130_fd_sc_hd__inv_2
X_2126_ _2127_/CLK _1808_/Y VGND VGND VPWR VPWR _1804_/A sky130_fd_sc_hd__dfxtp_4
X_2057_ _2137_/CLK DATA_FROM_HASH[6] VGND VGND VPWR VPWR _2057_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1008_ _1750_/A VGND VGND VPWR VPWR _1008_/X sky130_fd_sc_hd__buf_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1290_ _1892_/A _1279_/Y _1283_/X VGND VGND VPWR VPWR _1290_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_63_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1626_ _1585_/B _1624_/X _1681_/A VGND VGND VPWR VPWR _1628_/A sky130_fd_sc_hd__o21a_4
X_1557_ _2186_/Q _2187_/Q VGND VGND VPWR VPWR _1570_/C sky130_fd_sc_hd__nand2_4
XFILLER_39_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1488_ _1057_/A _1487_/Y _1057_/C _1389_/B VGND VGND VPWR VPWR _1488_/X sky130_fd_sc_hd__o22a_4
X_2109_ _2121_/CLK _1844_/Y VGND VGND VPWR VPWR _2109_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1273_ _1268_/Y _1269_/Y _1272_/X VGND VGND VPWR VPWR _1275_/A sky130_fd_sc_hd__a21o_4
X_1342_ _1342_/A VGND VGND VPWR VPWR _1342_/Y sky130_fd_sc_hd__inv_2
X_1411_ _2060_/Q VGND VGND VPWR VPWR _1412_/B sky130_fd_sc_hd__inv_2
XFILLER_51_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1609_ _1609_/A _1577_/A _1609_/C _1609_/D VGND VGND VPWR VPWR _1609_/X sky130_fd_sc_hd__and4_4
XFILLER_63_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1891_ _1042_/Y _1885_/X _1888_/X _1169_/Y _1890_/X VGND VGND VPWR VPWR _2090_/D
+ sky130_fd_sc_hd__o32ai_4
X_1960_ _1003_/A _1972_/C _1654_/A VGND VGND VPWR VPWR _1960_/X sky130_fd_sc_hd__a21o_4
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1256_ _1164_/X _2072_/Q _1166_/A VGND VGND VPWR VPWR _1256_/Y sky130_fd_sc_hd__a21oi_4
X_1325_ _1325_/A VGND VGND VPWR VPWR _1325_/X sky130_fd_sc_hd__buf_2
X_1187_ _1187_/A VGND VGND VPWR VPWR _1188_/A sky130_fd_sc_hd__inv_2
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_8_0_addressalyzerBlock.SPI_CLK clkbuf_4_9_0_addressalyzerBlock.SPI_CLK/A
+ VGND VGND VPWR VPWR _2216_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_3_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE2_1 _1883_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2090_ _2083_/CLK _2090_/D VGND VGND VPWR VPWR _2090_/Q sky130_fd_sc_hd__dfxtp_4
X_1110_ _1056_/Y VGND VGND VPWR VPWR _1298_/C sky130_fd_sc_hd__buf_2
XFILLER_61_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1041_ _1034_/Y _1036_/Y _1040_/X VGND VGND VPWR VPWR _1041_/Y sky130_fd_sc_hd__a21oi_4
X_1943_ _1943_/A VGND VGND VPWR VPWR _1944_/A sky130_fd_sc_hd__inv_2
X_1874_ _1874_/A _1867_/B _2039_/D VGND VGND VPWR VPWR _1874_/Y sky130_fd_sc_hd__nand3_4
XFILLER_56_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1239_ _1235_/Y _1238_/Y _1175_/X VGND VGND VPWR VPWR _1239_/Y sky130_fd_sc_hd__a21oi_4
X_1308_ _1449_/A VGND VGND VPWR VPWR _1436_/A sky130_fd_sc_hd__buf_2
XFILLER_64_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1590_ CLK_LED VGND VGND VPWR VPWR _1590_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2073_ _2137_/CLK _1931_/X VGND VGND VPWR VPWR _2073_/Q sky130_fd_sc_hd__dfxtp_4
X_2142_ _2142_/CLK _2142_/D VGND VGND VPWR VPWR _1175_/A sky130_fd_sc_hd__dfxtp_4
X_2211_ _2225_/CLK _2211_/D VGND VGND VPWR VPWR _1496_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1024_ _1024_/A _1016_/B VGND VGND VPWR VPWR _1024_/X sky130_fd_sc_hd__or2_4
XFILLER_34_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1788_ _1788_/A _1402_/Y _1803_/A _1787_/Y VGND VGND VPWR VPWR _1788_/Y sky130_fd_sc_hd__nor4_4
X_1926_ _1907_/Y _1909_/X _1905_/A _1712_/Y _1910_/X VGND VGND VPWR VPWR _1926_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1857_ _1922_/C _1857_/B _1857_/C VGND VGND VPWR VPWR _1857_/Y sky130_fd_sc_hd__nand3_4
XFILLER_57_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1711_ _1180_/B _2043_/Q _1188_/A VGND VGND VPWR VPWR _1711_/Y sky130_fd_sc_hd__o21ai_4
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1642_ _1582_/A _1647_/A _1661_/B VGND VGND VPWR VPWR _1642_/Y sky130_fd_sc_hd__nor3_4
XFILLER_6_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1573_ _1963_/A _1573_/B VGND VGND VPWR VPWR _2185_/D sky130_fd_sc_hd__nor2_4
X_2056_ _2056_/CLK DATA_FROM_HASH[5] VGND VGND VPWR VPWR _2048_/D sky130_fd_sc_hd__dfxtp_4
X_2125_ _2127_/CLK _2125_/D VGND VGND VPWR VPWR _1804_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_26_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1007_ _1504_/A VGND VGND VPWR VPWR _1750_/A sky130_fd_sc_hd__buf_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1909_ _1909_/A VGND VGND VPWR VPWR _1909_/X sky130_fd_sc_hd__buf_2
XFILLER_1_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1625_ _1504_/A VGND VGND VPWR VPWR _1681_/A sky130_fd_sc_hd__buf_2
X_1556_ _0997_/X _1545_/C _1555_/Y VGND VGND VPWR VPWR _2191_/D sky130_fd_sc_hd__o21a_4
XFILLER_39_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1487_ _1487_/A VGND VGND VPWR VPWR _1487_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2039_ _2016_/CLK _2039_/D VGND VGND VPWR VPWR _2039_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_52_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2108_ _2121_/CLK _1846_/Y VGND VGND VPWR VPWR _2108_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1410_ _1406_/X _1409_/Y _1175_/A VGND VGND VPWR VPWR _1414_/A sky130_fd_sc_hd__a21o_4
X_1272_ _1271_/Y _1272_/B VGND VGND VPWR VPWR _1272_/X sky130_fd_sc_hd__or2_4
X_1341_ _1338_/X _1339_/Y _1341_/C VGND VGND VPWR VPWR _1342_/A sky130_fd_sc_hd__nand3_4
XFILLER_36_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1608_ _1607_/X _1608_/B _1583_/Y VGND VGND VPWR VPWR _1609_/A sky130_fd_sc_hd__nor3_4
X_1539_ _2195_/Q _1525_/A _1538_/X VGND VGND VPWR VPWR _1539_/X sky130_fd_sc_hd__o21a_4
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1890_ _1889_/X VGND VGND VPWR VPWR _1890_/X sky130_fd_sc_hd__buf_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1255_ ID_toHost VGND VGND VPWR VPWR _1255_/Y sky130_fd_sc_hd__inv_2
X_1186_ _1189_/A _1186_/B VGND VGND VPWR VPWR _1187_/A sky130_fd_sc_hd__nor2_4
Xclkbuf_4_13_0_addressalyzerBlock.SPI_CLK clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/X
+ VGND VGND VPWR VPWR _2077_/CLK sky130_fd_sc_hd__clkbuf_1
X_1324_ _1315_/Y _1323_/Y _1040_/X VGND VGND VPWR VPWR _1324_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_64_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE2_2 _2094_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_7_0_m1_clk_local clkbuf_2_3_0_m1_clk_local/X VGND VGND VPWR VPWR _2121_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1040_ _1039_/X VGND VGND VPWR VPWR _1040_/X sky130_fd_sc_hd__buf_2
XFILLER_61_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1942_ _1419_/C _1863_/B _1886_/B _1737_/D VGND VGND VPWR VPWR _1943_/A sky130_fd_sc_hd__and4_4
XFILLER_21_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1873_ _1932_/A _1865_/X _1872_/Y VGND VGND VPWR VPWR _2096_/D sky130_fd_sc_hd__o21ai_4
XFILLER_9_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1238_ _1236_/Y _1170_/X _1237_/Y VGND VGND VPWR VPWR _1238_/Y sky130_fd_sc_hd__o21ai_4
X_1169_ _2090_/Q VGND VGND VPWR VPWR _1169_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1307_ _1307_/A _1307_/B _1306_/Y VGND VGND VPWR VPWR _2224_/D sky130_fd_sc_hd__and3_4
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2210_ _2216_/CLK _2210_/D VGND VGND VPWR VPWR _1499_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_53_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2141_ _2077_/CLK _1706_/Y VGND VGND VPWR VPWR _1172_/A sky130_fd_sc_hd__dfxtp_4
X_2072_ _2137_/CLK _1933_/X VGND VGND VPWR VPWR _2072_/Q sky130_fd_sc_hd__dfxtp_4
X_1023_ _1021_/Y _1003_/X _1022_/Y VGND VGND VPWR VPWR _1023_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_61_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1925_ _1904_/Y _1918_/A _1924_/Y VGND VGND VPWR VPWR _2076_/D sky130_fd_sc_hd__o21ai_4
XFILLER_34_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1787_ _1825_/A _1813_/C _1813_/D _1787_/D VGND VGND VPWR VPWR _1787_/Y sky130_fd_sc_hd__nand4_4
X_1856_ _1856_/A _1856_/B VGND VGND VPWR VPWR _2102_/D sky130_fd_sc_hd__xor2_4
XFILLER_40_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1572_ _2186_/Q _1571_/Y VGND VGND VPWR VPWR _1572_/Y sky130_fd_sc_hd__nor2_4
X_1710_ _1857_/C _1365_/A _1421_/Y VGND VGND VPWR VPWR _1731_/A sky130_fd_sc_hd__o21ai_4
X_1641_ _1582_/D VGND VGND VPWR VPWR _1661_/B sky130_fd_sc_hd__buf_2
X_2124_ _2127_/CLK _1810_/X VGND VGND VPWR VPWR _2124_/Q sky130_fd_sc_hd__dfxtp_4
X_1006_ _1863_/B VGND VGND VPWR VPWR _1504_/A sky130_fd_sc_hd__buf_2
X_2055_ _2216_/CLK DATA_FROM_HASH[4] VGND VGND VPWR VPWR _2055_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1839_ _1839_/A _1839_/B VGND VGND VPWR VPWR _2112_/D sky130_fd_sc_hd__xor2_4
X_1908_ _1907_/Y _1473_/B _1905_/X _1715_/Y _1889_/X VGND VGND VPWR VPWR _2083_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_22_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1624_ _1619_/Y _1621_/B _1577_/A _1585_/A VGND VGND VPWR VPWR _1624_/X sky130_fd_sc_hd__and4_4
X_1555_ _1554_/Y VGND VGND VPWR VPWR _1555_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2107_ _2110_/CLK _1848_/Y VGND VGND VPWR VPWR _1845_/A sky130_fd_sc_hd__dfxtp_4
X_1486_ _1486_/A VGND VGND VPWR VPWR _1498_/B sky130_fd_sc_hd__inv_2
XFILLER_54_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2038_ _2027_/CLK _2094_/Q VGND VGND VPWR VPWR _2032_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1340_ _1917_/A VGND VGND VPWR VPWR _1341_/C sky130_fd_sc_hd__buf_2
XFILLER_5_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1271_ _1772_/A _1365_/A VGND VGND VPWR VPWR _1271_/Y sky130_fd_sc_hd__nor2_4
XFILLER_36_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1469_ _1189_/A _1191_/A _1723_/A _2047_/Q VGND VGND VPWR VPWR _1469_/Y sky130_fd_sc_hd__a2bb2oi_4
X_1607_ _1575_/Y VGND VGND VPWR VPWR _1607_/X sky130_fd_sc_hd__buf_2
X_1538_ _2196_/Q _1526_/A _1535_/X VGND VGND VPWR VPWR _1538_/X sky130_fd_sc_hd__o21a_4
XFILLER_63_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1323_ _1317_/Y _1318_/X _1323_/C VGND VGND VPWR VPWR _1323_/Y sky130_fd_sc_hd__nand3_4
XFILLER_64_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1254_ _1159_/X _1490_/A _1161_/X VGND VGND VPWR VPWR _1254_/Y sky130_fd_sc_hd__a21oi_4
X_1185_ _1185_/A VGND VGND VPWR VPWR _1186_/B sky130_fd_sc_hd__inv_2
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE2_3 _2085_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1941_ _1935_/A _1753_/A _2067_/Q _1185_/A _1940_/Y VGND VGND VPWR VPWR _1941_/X
+ sky130_fd_sc_hd__a32o_4
X_1872_ _1874_/A _1867_/B _1872_/C VGND VGND VPWR VPWR _1872_/Y sky130_fd_sc_hd__nand3_4
XFILLER_14_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1306_ _1283_/X _1086_/X VGND VGND VPWR VPWR _1306_/Y sky130_fd_sc_hd__nand2_4
XFILLER_64_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1168_ _1163_/Y _1159_/X _1167_/Y VGND VGND VPWR VPWR _1168_/Y sky130_fd_sc_hd__o21ai_4
X_1237_ _1171_/X _2097_/Q _1172_/A VGND VGND VPWR VPWR _1237_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_37_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1099_ _1070_/X _1097_/Y _1446_/A VGND VGND VPWR VPWR _1099_/X sky130_fd_sc_hd__a21o_4
XFILLER_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2140_ _2069_/CLK _2140_/D VGND VGND VPWR VPWR _1347_/A sky130_fd_sc_hd__dfxtp_4
X_2071_ _2056_/CLK _1936_/Y VGND VGND VPWR VPWR _1462_/A sky130_fd_sc_hd__dfxtp_4
X_1022_ _2219_/Q _1004_/X _1008_/X VGND VGND VPWR VPWR _1022_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_61_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1924_ _1924_/A _1918_/B _2076_/Q VGND VGND VPWR VPWR _1924_/Y sky130_fd_sc_hd__nand3_4
X_1855_ _2103_/Q _1854_/Y VGND VGND VPWR VPWR _1855_/X sky130_fd_sc_hd__xor2_4
X_1786_ _1785_/Y VGND VGND VPWR VPWR _1787_/D sky130_fd_sc_hd__inv_2
XFILLER_52_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1571_ SPI_CLK_RESET_N VGND VGND VPWR VPWR _1571_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1640_ _1607_/X _1646_/C _1639_/Y VGND VGND VPWR VPWR _1640_/Y sky130_fd_sc_hd__a21oi_4
X_2123_ _2127_/CLK _2123_/D VGND VGND VPWR VPWR _1769_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_26_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1005_ _2004_/Q VGND VGND VPWR VPWR _1863_/B sky130_fd_sc_hd__inv_2
X_2054_ _2216_/CLK DATA_FROM_HASH[3] VGND VGND VPWR VPWR _2054_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1838_ _1838_/A _1838_/B VGND VGND VPWR VPWR _1839_/B sky130_fd_sc_hd__nor2_4
X_1907_ _1907_/A VGND VGND VPWR VPWR _1907_/Y sky130_fd_sc_hd__inv_2
X_1769_ _1769_/A VGND VGND VPWR VPWR _1803_/A sky130_fd_sc_hd__inv_2
XFILLER_45_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1485_ _1097_/Y _1490_/A _1482_/Y _1483_/X _1484_/X VGND VGND VPWR VPWR _1486_/A
+ sky130_fd_sc_hd__a2111o_4
X_1623_ _1609_/C _1621_/X _1622_/Y VGND VGND VPWR VPWR _2178_/D sky130_fd_sc_hd__o21a_4
X_1554_ _1549_/A _1535_/X _1553_/Y VGND VGND VPWR VPWR _1554_/Y sky130_fd_sc_hd__nand3_4
.ends

