VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO decred_top
  CLASS BLOCK ;
  FOREIGN decred_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 3400.000 ;
  PIN CLK_LED
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1370.920 4.000 1371.520 ;
    END
  END CLK_LED
  PIN EXT_RESET_N_fromHost
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2778.490 0.000 2778.770 4.000 ;
    END
  END EXT_RESET_N_fromHost
  PIN EXT_RESET_N_toClient
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 464.690 0.000 464.970 4.000 ;
    END
  END EXT_RESET_N_toClient
  PIN HASH_LED
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END HASH_LED
  PIN ID_fromClient
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2739.080 4.000 2739.680 ;
    END
  END ID_fromClient
  PIN ID_toHost
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2796.000 2027.800 2800.000 2028.400 ;
    END
  END ID_toHost
  PIN IRQ_OUT_fromClient
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2796.890 3396.000 2797.170 3400.000 ;
    END
  END IRQ_OUT_fromClient
  PIN IRQ_OUT_toHost
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1390.210 0.000 1390.490 4.000 ;
    END
  END IRQ_OUT_toHost
  PIN M1_CLK_IN
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1852.970 0.000 1853.250 4.000 ;
    END
  END M1_CLK_IN
  PIN M1_CLK_SELECT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1409.530 3396.000 1409.810 3400.000 ;
    END
  END M1_CLK_SELECT
  PIN MISO_fromClient
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2796.000 659.640 2800.000 660.240 ;
    END
  END MISO_fromClient
  PIN MISO_toHost
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END MISO_toHost
  PIN MOSI_fromHost
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2335.050 3396.000 2335.330 3400.000 ;
    END
  END MOSI_fromHost
  PIN MOSI_toClient
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2796.000 2711.880 2800.000 2712.480 ;
    END
  END MOSI_toClient
  PIN PLL_INPUT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1872.290 3396.000 1872.570 3400.000 ;
    END
  END PLL_INPUT
  PIN S1_CLK_IN
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 4.000 ;
    END
  END S1_CLK_IN
  PIN S1_CLK_SELECT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.250 3396.000 21.530 3400.000 ;
    END
  END S1_CLK_SELECT
  PIN SCLK_fromHost
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 946.770 3396.000 947.050 3400.000 ;
    END
  END SCLK_fromHost
  PIN SCLK_toClient
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2055.000 4.000 2055.600 ;
    END
  END SCLK_toClient
  PIN SCSN_fromHost
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2315.730 0.000 2316.010 4.000 ;
    END
  END SCSN_fromHost
  PIN SCSN_toClient
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 484.010 3396.000 484.290 3400.000 ;
    END
  END SCSN_toClient
  PIN SPI_CLK_RESET_N
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1343.720 2800.000 1344.320 ;
    END
  END SPI_CLK_RESET_N
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 36.240 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 36.240 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2794.040 3389.205 ;
      LAYER met1 ;
        RECT 2.830 10.640 2797.190 3389.360 ;
      LAYER met2 ;
        RECT 2.860 3395.720 20.970 3396.000 ;
        RECT 21.810 3395.720 483.730 3396.000 ;
        RECT 484.570 3395.720 946.490 3396.000 ;
        RECT 947.330 3395.720 1409.250 3396.000 ;
        RECT 1410.090 3395.720 1872.010 3396.000 ;
        RECT 1872.850 3395.720 2334.770 3396.000 ;
        RECT 2335.610 3395.720 2796.610 3396.000 ;
        RECT 2.860 4.280 2797.160 3395.720 ;
        RECT 3.410 4.000 464.410 4.280 ;
        RECT 465.250 4.000 927.170 4.280 ;
        RECT 928.010 4.000 1389.930 4.280 ;
        RECT 1390.770 4.000 1852.690 4.280 ;
        RECT 1853.530 4.000 2315.450 4.280 ;
        RECT 2316.290 4.000 2778.210 4.280 ;
        RECT 2779.050 4.000 2797.160 4.280 ;
      LAYER met3 ;
        RECT 4.000 2740.080 2796.000 3389.285 ;
        RECT 4.400 2738.680 2796.000 2740.080 ;
        RECT 4.000 2712.880 2796.000 2738.680 ;
        RECT 4.000 2711.480 2795.600 2712.880 ;
        RECT 4.000 2056.000 2796.000 2711.480 ;
        RECT 4.400 2054.600 2796.000 2056.000 ;
        RECT 4.000 2028.800 2796.000 2054.600 ;
        RECT 4.000 2027.400 2795.600 2028.800 ;
        RECT 4.000 1371.920 2796.000 2027.400 ;
        RECT 4.400 1370.520 2796.000 1371.920 ;
        RECT 4.000 1344.720 2796.000 1370.520 ;
        RECT 4.000 1343.320 2795.600 1344.720 ;
        RECT 4.000 687.840 2796.000 1343.320 ;
        RECT 4.400 686.440 2796.000 687.840 ;
        RECT 4.000 660.640 2796.000 686.440 ;
        RECT 4.000 659.240 2795.600 660.640 ;
        RECT 4.000 10.715 2796.000 659.240 ;
      LAYER met4 ;
        RECT 21.040 36.640 2787.440 3389.360 ;
        RECT 21.040 10.640 327.840 36.640 ;
        RECT 330.240 10.640 404.640 36.640 ;
        RECT 407.040 10.640 2787.440 36.640 ;
      LAYER met5 ;
        RECT 1132.180 506.300 1145.740 507.900 ;
  END
END decred_top
END LIBRARY

