VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO decred_controller
  CLASS BLOCK ;
  FOREIGN decred_controller ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN CLK_LED
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END CLK_LED
  PIN DATA_AVAILABLE[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 95.770 196.000 96.050 200.000 ;
    END
  END DATA_AVAILABLE[0]
  PIN DATA_AVAILABLE[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 196.000 74.890 200.000 ;
    END
  END DATA_AVAILABLE[1]
  PIN DATA_AVAILABLE[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END DATA_AVAILABLE[2]
  PIN DATA_AVAILABLE[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 159.250 196.000 159.530 200.000 ;
    END
  END DATA_AVAILABLE[3]
  PIN DATA_AVAILABLE[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END DATA_AVAILABLE[4]
  PIN DATA_FROM_HASH[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END DATA_FROM_HASH[0]
  PIN DATA_FROM_HASH[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 138.090 196.000 138.370 200.000 ;
    END
  END DATA_FROM_HASH[1]
  PIN DATA_FROM_HASH[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.130 196.000 11.410 200.000 ;
    END
  END DATA_FROM_HASH[2]
  PIN DATA_FROM_HASH[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END DATA_FROM_HASH[3]
  PIN DATA_FROM_HASH[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 61.240 200.000 61.840 ;
    END
  END DATA_FROM_HASH[4]
  PIN DATA_FROM_HASH[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.570 196.000 63.850 200.000 ;
    END
  END DATA_FROM_HASH[5]
  PIN DATA_FROM_HASH[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END DATA_FROM_HASH[6]
  PIN DATA_FROM_HASH[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END DATA_FROM_HASH[7]
  PIN DATA_TO_HASH[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 170.290 196.000 170.570 200.000 ;
    END
  END DATA_TO_HASH[0]
  PIN DATA_TO_HASH[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END DATA_TO_HASH[1]
  PIN DATA_TO_HASH[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END DATA_TO_HASH[2]
  PIN DATA_TO_HASH[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 21.250 196.000 21.530 200.000 ;
    END
  END DATA_TO_HASH[3]
  PIN DATA_TO_HASH[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 15.000 200.000 15.600 ;
    END
  END DATA_TO_HASH[4]
  PIN DATA_TO_HASH[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 108.840 200.000 109.440 ;
    END
  END DATA_TO_HASH[5]
  PIN DATA_TO_HASH[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END DATA_TO_HASH[6]
  PIN DATA_TO_HASH[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 105.890 196.000 106.170 200.000 ;
    END
  END DATA_TO_HASH[7]
  PIN EXT_RESET_N_fromHost
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END EXT_RESET_N_fromHost
  PIN EXT_RESET_N_toClient
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END EXT_RESET_N_toClient
  PIN HASH_ADDR[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 149.130 196.000 149.410 200.000 ;
    END
  END HASH_ADDR[0]
  PIN HASH_ADDR[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END HASH_ADDR[1]
  PIN HASH_ADDR[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.050 196.000 127.330 200.000 ;
    END
  END HASH_ADDR[2]
  PIN HASH_ADDR[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END HASH_ADDR[3]
  PIN HASH_ADDR[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END HASH_ADDR[4]
  PIN HASH_ADDR[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 53.450 196.000 53.730 200.000 ;
    END
  END HASH_ADDR[5]
  PIN HASH_EN
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END HASH_EN
  PIN HASH_LED
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 77.560 200.000 78.160 ;
    END
  END HASH_LED
  PIN ID_fromClient
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END ID_fromClient
  PIN ID_toHost
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 125.160 200.000 125.760 ;
    END
  END ID_toHost
  PIN IRQ_OUT_fromClient
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END IRQ_OUT_fromClient
  PIN IRQ_OUT_toHost
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END IRQ_OUT_toHost
  PIN M1_CLK_IN
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END M1_CLK_IN
  PIN M1_CLK_SELECT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END M1_CLK_SELECT
  PIN MACRO_RD_SELECT[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END MACRO_RD_SELECT[0]
  PIN MACRO_RD_SELECT[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END MACRO_RD_SELECT[1]
  PIN MACRO_RD_SELECT[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END MACRO_RD_SELECT[2]
  PIN MACRO_RD_SELECT[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 32.290 196.000 32.570 200.000 ;
    END
  END MACRO_RD_SELECT[3]
  PIN MACRO_RD_SELECT[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END MACRO_RD_SELECT[4]
  PIN MACRO_WR_SELECT[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 180.410 196.000 180.690 200.000 ;
    END
  END MACRO_WR_SELECT[0]
  PIN MACRO_WR_SELECT[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 46.280 200.000 46.880 ;
    END
  END MACRO_WR_SELECT[1]
  PIN MACRO_WR_SELECT[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END MACRO_WR_SELECT[2]
  PIN MACRO_WR_SELECT[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.930 196.000 117.210 200.000 ;
    END
  END MACRO_WR_SELECT[3]
  PIN MACRO_WR_SELECT[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 191.450 196.000 191.730 200.000 ;
    END
  END MACRO_WR_SELECT[4]
  PIN MISO_fromClient
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 92.520 200.000 93.120 ;
    END
  END MISO_fromClient
  PIN MISO_toHost
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 29.960 200.000 30.560 ;
    END
  END MISO_toHost
  PIN MOSI_fromHost
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END MOSI_fromHost
  PIN MOSI_toClient
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 187.720 200.000 188.320 ;
    END
  END MOSI_toClient
  PIN PLL_INPUT
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 171.400 200.000 172.000 ;
    END
  END PLL_INPUT
  PIN S1_CLK_IN
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END S1_CLK_IN
  PIN S1_CLK_SELECT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 84.730 196.000 85.010 200.000 ;
    END
  END S1_CLK_SELECT
  PIN SCLK_fromHost
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 156.440 200.000 157.040 ;
    END
  END SCLK_fromHost
  PIN SCLK_toClient
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END SCLK_toClient
  PIN SCSN_fromHost
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 140.120 200.000 140.720 ;
    END
  END SCSN_fromHost
  PIN SCSN_toClient
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END SCSN_toClient
  PIN SPI_CLK_RESET_N
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.410 196.000 42.690 200.000 ;
    END
  END SPI_CLK_RESET_N
  PIN m1_clk_local
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END m1_clk_local
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.895 187.765 ;
      LAYER met1 ;
        RECT 2.830 9.560 194.970 188.320 ;
      LAYER met2 ;
        RECT 2.860 195.720 10.850 196.000 ;
        RECT 11.690 195.720 20.970 196.000 ;
        RECT 21.810 195.720 32.010 196.000 ;
        RECT 32.850 195.720 42.130 196.000 ;
        RECT 42.970 195.720 53.170 196.000 ;
        RECT 54.010 195.720 63.290 196.000 ;
        RECT 64.130 195.720 74.330 196.000 ;
        RECT 75.170 195.720 84.450 196.000 ;
        RECT 85.290 195.720 95.490 196.000 ;
        RECT 96.330 195.720 105.610 196.000 ;
        RECT 106.450 195.720 116.650 196.000 ;
        RECT 117.490 195.720 126.770 196.000 ;
        RECT 127.610 195.720 137.810 196.000 ;
        RECT 138.650 195.720 148.850 196.000 ;
        RECT 149.690 195.720 158.970 196.000 ;
        RECT 159.810 195.720 170.010 196.000 ;
        RECT 170.850 195.720 180.130 196.000 ;
        RECT 180.970 195.720 191.170 196.000 ;
        RECT 192.010 195.720 194.950 196.000 ;
        RECT 2.860 4.280 194.950 195.720 ;
        RECT 3.410 4.000 12.690 4.280 ;
        RECT 13.530 4.000 23.730 4.280 ;
        RECT 24.570 4.000 33.850 4.280 ;
        RECT 34.690 4.000 44.890 4.280 ;
        RECT 45.730 4.000 55.010 4.280 ;
        RECT 55.850 4.000 66.050 4.280 ;
        RECT 66.890 4.000 76.170 4.280 ;
        RECT 77.010 4.000 87.210 4.280 ;
        RECT 88.050 4.000 97.330 4.280 ;
        RECT 98.170 4.000 108.370 4.280 ;
        RECT 109.210 4.000 118.490 4.280 ;
        RECT 119.330 4.000 129.530 4.280 ;
        RECT 130.370 4.000 140.570 4.280 ;
        RECT 141.410 4.000 150.690 4.280 ;
        RECT 151.530 4.000 161.730 4.280 ;
        RECT 162.570 4.000 171.850 4.280 ;
        RECT 172.690 4.000 182.890 4.280 ;
        RECT 183.730 4.000 193.010 4.280 ;
        RECT 193.850 4.000 194.950 4.280 ;
      LAYER met3 ;
        RECT 4.400 191.400 196.000 192.265 ;
        RECT 4.000 188.720 196.000 191.400 ;
        RECT 4.000 187.320 195.600 188.720 ;
        RECT 4.000 176.480 196.000 187.320 ;
        RECT 4.400 175.080 196.000 176.480 ;
        RECT 4.000 172.400 196.000 175.080 ;
        RECT 4.000 171.000 195.600 172.400 ;
        RECT 4.000 161.520 196.000 171.000 ;
        RECT 4.400 160.120 196.000 161.520 ;
        RECT 4.000 157.440 196.000 160.120 ;
        RECT 4.000 156.040 195.600 157.440 ;
        RECT 4.000 145.200 196.000 156.040 ;
        RECT 4.400 143.800 196.000 145.200 ;
        RECT 4.000 141.120 196.000 143.800 ;
        RECT 4.000 139.720 195.600 141.120 ;
        RECT 4.000 130.240 196.000 139.720 ;
        RECT 4.400 128.840 196.000 130.240 ;
        RECT 4.000 126.160 196.000 128.840 ;
        RECT 4.000 124.760 195.600 126.160 ;
        RECT 4.000 113.920 196.000 124.760 ;
        RECT 4.400 112.520 196.000 113.920 ;
        RECT 4.000 109.840 196.000 112.520 ;
        RECT 4.000 108.440 195.600 109.840 ;
        RECT 4.000 98.960 196.000 108.440 ;
        RECT 4.400 97.560 196.000 98.960 ;
        RECT 4.000 93.520 196.000 97.560 ;
        RECT 4.000 92.120 195.600 93.520 ;
        RECT 4.000 82.640 196.000 92.120 ;
        RECT 4.400 81.240 196.000 82.640 ;
        RECT 4.000 78.560 196.000 81.240 ;
        RECT 4.000 77.160 195.600 78.560 ;
        RECT 4.000 67.680 196.000 77.160 ;
        RECT 4.400 66.280 196.000 67.680 ;
        RECT 4.000 62.240 196.000 66.280 ;
        RECT 4.000 60.840 195.600 62.240 ;
        RECT 4.000 51.360 196.000 60.840 ;
        RECT 4.400 49.960 196.000 51.360 ;
        RECT 4.000 47.280 196.000 49.960 ;
        RECT 4.000 45.880 195.600 47.280 ;
        RECT 4.000 36.400 196.000 45.880 ;
        RECT 4.400 35.000 196.000 36.400 ;
        RECT 4.000 30.960 196.000 35.000 ;
        RECT 4.000 29.560 195.600 30.960 ;
        RECT 4.000 20.080 196.000 29.560 ;
        RECT 4.400 18.680 196.000 20.080 ;
        RECT 4.000 16.000 196.000 18.680 ;
        RECT 4.000 14.600 195.600 16.000 ;
        RECT 4.000 10.715 196.000 14.600 ;
      LAYER met4 ;
        RECT 62.855 10.640 97.440 187.920 ;
        RECT 99.840 10.640 176.240 187.920 ;
  END
END decred_controller
END LIBRARY

