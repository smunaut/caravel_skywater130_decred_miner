magic
tech sky130A
magscale 1 2
timestamp 1608049295
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 566 2128 38824 37584
<< metal2 >>
rect 2778 39200 2834 40000
rect 5170 39200 5226 40000
rect 7562 39200 7618 40000
rect 9770 39200 9826 40000
rect 12162 39200 12218 40000
rect 14554 39200 14610 40000
rect 16946 39200 17002 40000
rect 19338 39200 19394 40000
rect 21546 39200 21602 40000
rect 23938 39200 23994 40000
rect 26330 39200 26386 40000
rect 28722 39200 28778 40000
rect 31114 39200 31170 40000
rect 33322 39200 33378 40000
rect 35714 39200 35770 40000
rect 38106 39200 38162 40000
rect 570 0 626 800
rect 2778 0 2834 800
rect 5170 0 5226 800
rect 7562 0 7618 800
rect 9954 0 10010 800
rect 12346 0 12402 800
rect 14554 0 14610 800
rect 16946 0 17002 800
rect 19338 0 19394 800
rect 21730 0 21786 800
rect 24122 0 24178 800
rect 26330 0 26386 800
rect 28722 0 28778 800
rect 31114 0 31170 800
rect 33506 0 33562 800
rect 35898 0 35954 800
rect 38106 0 38162 800
<< obsm2 >>
rect 572 39144 2722 39200
rect 2890 39144 5114 39200
rect 5282 39144 7506 39200
rect 7674 39144 9714 39200
rect 9882 39144 12106 39200
rect 12274 39144 14498 39200
rect 14666 39144 16890 39200
rect 17058 39144 19282 39200
rect 19450 39144 21490 39200
rect 21658 39144 23882 39200
rect 24050 39144 26274 39200
rect 26442 39144 28666 39200
rect 28834 39144 31058 39200
rect 31226 39144 33266 39200
rect 33434 39144 35658 39200
rect 35826 39144 38050 39200
rect 572 856 38160 39144
rect 682 800 2722 856
rect 2890 800 5114 856
rect 5282 800 7506 856
rect 7674 800 9898 856
rect 10066 800 12290 856
rect 12458 800 14498 856
rect 14666 800 16890 856
rect 17058 800 19282 856
rect 19450 800 21674 856
rect 21842 800 24066 856
rect 24234 800 26274 856
rect 26442 800 28666 856
rect 28834 800 31058 856
rect 31226 800 33450 856
rect 33618 800 35842 856
rect 36010 800 38050 856
<< metal3 >>
rect 0 38904 800 39024
rect 39200 37272 40000 37392
rect 0 35368 800 35488
rect 39200 33736 40000 33856
rect 0 32104 800 32224
rect 39200 30472 40000 30592
rect 0 28568 800 28688
rect 39200 26936 40000 27056
rect 0 25032 800 25152
rect 39200 23400 40000 23520
rect 0 21496 800 21616
rect 39200 19864 40000 19984
rect 0 17960 800 18080
rect 39200 16328 40000 16448
rect 0 14696 800 14816
rect 39200 13064 40000 13184
rect 0 11160 800 11280
rect 39200 9528 40000 9648
rect 0 7624 800 7744
rect 39200 5992 40000 6112
rect 0 4088 800 4208
rect 39200 2456 40000 2576
<< obsm3 >>
rect 880 38824 39200 38997
rect 800 37472 39200 38824
rect 800 37192 39120 37472
rect 800 35568 39200 37192
rect 880 35288 39200 35568
rect 800 33936 39200 35288
rect 800 33656 39120 33936
rect 800 32304 39200 33656
rect 880 32024 39200 32304
rect 800 30672 39200 32024
rect 800 30392 39120 30672
rect 800 28768 39200 30392
rect 880 28488 39200 28768
rect 800 27136 39200 28488
rect 800 26856 39120 27136
rect 800 25232 39200 26856
rect 880 24952 39200 25232
rect 800 23600 39200 24952
rect 800 23320 39120 23600
rect 800 21696 39200 23320
rect 880 21416 39200 21696
rect 800 20064 39200 21416
rect 800 19784 39120 20064
rect 800 18160 39200 19784
rect 880 17880 39200 18160
rect 800 16528 39200 17880
rect 800 16248 39120 16528
rect 800 14896 39200 16248
rect 880 14616 39200 14896
rect 800 13264 39200 14616
rect 800 12984 39120 13264
rect 800 11360 39200 12984
rect 880 11080 39200 11360
rect 800 9728 39200 11080
rect 800 9448 39120 9728
rect 800 7824 39200 9448
rect 880 7544 39200 7824
rect 800 6192 39200 7544
rect 800 5912 39120 6192
rect 800 4288 39200 5912
rect 880 4008 39200 4288
rect 800 2656 39200 4008
rect 800 2376 39120 2656
rect 800 2143 39200 2376
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
<< obsm4 >>
rect 18643 2128 19488 37584
rect 19968 2128 35248 37584
<< labels >>
rlabel metal3 s 0 21496 800 21616 6 CLK_LED
port 1 nsew default output
rlabel metal2 s 9770 39200 9826 40000 6 DATA_AVAILABLE
port 2 nsew default input
rlabel metal2 s 5170 39200 5226 40000 6 DATA_FROM_HASH[0]
port 3 nsew default input
rlabel metal3 s 0 35368 800 35488 6 DATA_FROM_HASH[1]
port 4 nsew default input
rlabel metal2 s 23938 39200 23994 40000 6 DATA_FROM_HASH[2]
port 5 nsew default input
rlabel metal2 s 21730 0 21786 800 6 DATA_FROM_HASH[3]
port 6 nsew default input
rlabel metal2 s 26330 0 26386 800 6 DATA_FROM_HASH[4]
port 7 nsew default input
rlabel metal2 s 19338 39200 19394 40000 6 DATA_FROM_HASH[5]
port 8 nsew default input
rlabel metal3 s 0 25032 800 25152 6 DATA_FROM_HASH[6]
port 9 nsew default input
rlabel metal3 s 39200 37272 40000 37392 6 DATA_FROM_HASH[7]
port 10 nsew default input
rlabel metal3 s 39200 19864 40000 19984 6 DATA_TO_HASH[0]
port 11 nsew default output
rlabel metal2 s 2778 39200 2834 40000 6 DATA_TO_HASH[1]
port 12 nsew default output
rlabel metal2 s 28722 0 28778 800 6 DATA_TO_HASH[2]
port 13 nsew default output
rlabel metal3 s 0 4088 800 4208 6 DATA_TO_HASH[3]
port 14 nsew default output
rlabel metal2 s 26330 39200 26386 40000 6 DATA_TO_HASH[4]
port 15 nsew default output
rlabel metal2 s 5170 0 5226 800 6 DATA_TO_HASH[5]
port 16 nsew default output
rlabel metal3 s 39200 2456 40000 2576 6 DATA_TO_HASH[6]
port 17 nsew default output
rlabel metal3 s 0 28568 800 28688 6 DATA_TO_HASH[7]
port 18 nsew default output
rlabel metal3 s 39200 9528 40000 9648 6 EXT_RESET_N_fromHost
port 19 nsew default input
rlabel metal3 s 39200 30472 40000 30592 6 EXT_RESET_N_toClient
port 20 nsew default output
rlabel metal2 s 38106 0 38162 800 6 HASH_ADDR[0]
port 21 nsew default output
rlabel metal2 s 12162 39200 12218 40000 6 HASH_ADDR[1]
port 22 nsew default output
rlabel metal3 s 0 7624 800 7744 6 HASH_ADDR[2]
port 23 nsew default output
rlabel metal2 s 35898 0 35954 800 6 HASH_ADDR[3]
port 24 nsew default output
rlabel metal2 s 21546 39200 21602 40000 6 HASH_ADDR[4]
port 25 nsew default output
rlabel metal2 s 12346 0 12402 800 6 HASH_ADDR[5]
port 26 nsew default output
rlabel metal2 s 16946 39200 17002 40000 6 HASH_EN
port 27 nsew default output
rlabel metal2 s 33506 0 33562 800 6 HASH_LED
port 28 nsew default output
rlabel metal2 s 38106 39200 38162 40000 6 ID_fromClient
port 29 nsew default input
rlabel metal3 s 0 38904 800 39024 6 ID_toHost
port 30 nsew default output
rlabel metal2 s 16946 0 17002 800 6 IRQ_OUT_fromClient
port 31 nsew default input
rlabel metal3 s 39200 23400 40000 23520 6 IRQ_OUT_toHost
port 32 nsew default output
rlabel metal3 s 0 11160 800 11280 6 M1_CLK_IN
port 33 nsew default input
rlabel metal3 s 39200 33736 40000 33856 6 M1_CLK_SELECT
port 34 nsew default input
rlabel metal3 s 39200 5992 40000 6112 6 MACRO_RD_SELECT
port 35 nsew default output
rlabel metal2 s 9954 0 10010 800 6 MACRO_WR_SELECT
port 36 nsew default output
rlabel metal2 s 7562 0 7618 800 6 MISO_fromClient
port 37 nsew default input
rlabel metal2 s 31114 0 31170 800 6 MISO_toHost
port 38 nsew default output
rlabel metal2 s 24122 0 24178 800 6 MOSI_fromHost
port 39 nsew default input
rlabel metal2 s 19338 0 19394 800 6 MOSI_toClient
port 40 nsew default output
rlabel metal2 s 14554 0 14610 800 6 PLL_INPUT
port 41 nsew default input
rlabel metal3 s 0 32104 800 32224 6 S1_CLK_IN
port 42 nsew default input
rlabel metal2 s 2778 0 2834 800 6 S1_CLK_SELECT
port 43 nsew default input
rlabel metal2 s 28722 39200 28778 40000 6 SCLK_fromHost
port 44 nsew default input
rlabel metal3 s 39200 16328 40000 16448 6 SCLK_toClient
port 45 nsew default output
rlabel metal3 s 0 17960 800 18080 6 SCSN_fromHost
port 46 nsew default input
rlabel metal2 s 14554 39200 14610 40000 6 SCSN_toClient
port 47 nsew default output
rlabel metal2 s 31114 39200 31170 40000 6 SPI_CLK_RESET_N
port 48 nsew default input
rlabel metal3 s 39200 26936 40000 27056 6 THREAD_COUNT[0]
port 49 nsew default input
rlabel metal3 s 39200 13064 40000 13184 6 THREAD_COUNT[1]
port 50 nsew default input
rlabel metal2 s 570 0 626 800 6 THREAD_COUNT[2]
port 51 nsew default input
rlabel metal2 s 33322 39200 33378 40000 6 THREAD_COUNT[3]
port 52 nsew default input
rlabel metal2 s 35714 39200 35770 40000 6 m1_clk_local
port 53 nsew default output
rlabel metal3 s 0 14696 800 14816 6 one
port 54 nsew default output
rlabel metal2 s 7562 39200 7618 40000 6 zero
port 55 nsew default output
rlabel metal4 s 4208 2128 4528 37584 6 VPWR
port 56 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 VGND
port 57 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 40000 40000
string LEFview TRUE
<< end >>
