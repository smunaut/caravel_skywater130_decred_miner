VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO decred_controller
  CLASS BLOCK ;
  FOREIGN decred_controller ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN CLK_LED
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END CLK_LED
  PIN DATA_AVAILABLE
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 196.000 49.130 200.000 ;
    END
  END DATA_AVAILABLE
  PIN DATA_FROM_HASH[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.850 196.000 26.130 200.000 ;
    END
  END DATA_FROM_HASH[0]
  PIN DATA_FROM_HASH[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END DATA_FROM_HASH[1]
  PIN DATA_FROM_HASH[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 119.690 196.000 119.970 200.000 ;
    END
  END DATA_FROM_HASH[2]
  PIN DATA_FROM_HASH[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END DATA_FROM_HASH[3]
  PIN DATA_FROM_HASH[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END DATA_FROM_HASH[4]
  PIN DATA_FROM_HASH[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.690 196.000 96.970 200.000 ;
    END
  END DATA_FROM_HASH[5]
  PIN DATA_FROM_HASH[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END DATA_FROM_HASH[6]
  PIN DATA_FROM_HASH[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 186.360 200.000 186.960 ;
    END
  END DATA_FROM_HASH[7]
  PIN DATA_TO_HASH[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 99.320 200.000 99.920 ;
    END
  END DATA_TO_HASH[0]
  PIN DATA_TO_HASH[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 13.890 196.000 14.170 200.000 ;
    END
  END DATA_TO_HASH[1]
  PIN DATA_TO_HASH[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END DATA_TO_HASH[2]
  PIN DATA_TO_HASH[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END DATA_TO_HASH[3]
  PIN DATA_TO_HASH[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 131.650 196.000 131.930 200.000 ;
    END
  END DATA_TO_HASH[4]
  PIN DATA_TO_HASH[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END DATA_TO_HASH[5]
  PIN DATA_TO_HASH[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 12.280 200.000 12.880 ;
    END
  END DATA_TO_HASH[6]
  PIN DATA_TO_HASH[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END DATA_TO_HASH[7]
  PIN EXT_RESET_N_fromHost
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 47.640 200.000 48.240 ;
    END
  END EXT_RESET_N_fromHost
  PIN EXT_RESET_N_toClient
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 152.360 200.000 152.960 ;
    END
  END EXT_RESET_N_toClient
  PIN HASH_ADDR[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END HASH_ADDR[0]
  PIN HASH_ADDR[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 60.810 196.000 61.090 200.000 ;
    END
  END HASH_ADDR[1]
  PIN HASH_ADDR[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END HASH_ADDR[2]
  PIN HASH_ADDR[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END HASH_ADDR[3]
  PIN HASH_ADDR[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.730 196.000 108.010 200.000 ;
    END
  END HASH_ADDR[4]
  PIN HASH_ADDR[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END HASH_ADDR[5]
  PIN HASH_EN
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 84.730 196.000 85.010 200.000 ;
    END
  END HASH_EN
  PIN HASH_LED
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END HASH_LED
  PIN ID_fromClient
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 190.530 196.000 190.810 200.000 ;
    END
  END ID_fromClient
  PIN ID_toHost
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END ID_toHost
  PIN IRQ_OUT_fromClient
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END IRQ_OUT_fromClient
  PIN IRQ_OUT_toHost
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 117.000 200.000 117.600 ;
    END
  END IRQ_OUT_toHost
  PIN M1_CLK_IN
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END M1_CLK_IN
  PIN M1_CLK_SELECT
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 168.680 200.000 169.280 ;
    END
  END M1_CLK_SELECT
  PIN MACRO_RD_SELECT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 29.960 200.000 30.560 ;
    END
  END MACRO_RD_SELECT
  PIN MACRO_WR_SELECT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END MACRO_WR_SELECT
  PIN MISO_fromClient
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END MISO_fromClient
  PIN MISO_toHost
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END MISO_toHost
  PIN MOSI_fromHost
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END MOSI_fromHost
  PIN MOSI_toClient
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END MOSI_toClient
  PIN PLL_INPUT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END PLL_INPUT
  PIN S1_CLK_IN
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END S1_CLK_IN
  PIN S1_CLK_SELECT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END S1_CLK_SELECT
  PIN SCLK_fromHost
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 143.610 196.000 143.890 200.000 ;
    END
  END SCLK_fromHost
  PIN SCLK_toClient
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 81.640 200.000 82.240 ;
    END
  END SCLK_toClient
  PIN SCSN_fromHost
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END SCSN_fromHost
  PIN SCSN_toClient
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.770 196.000 73.050 200.000 ;
    END
  END SCSN_toClient
  PIN SPI_CLK_RESET_N
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 155.570 196.000 155.850 200.000 ;
    END
  END SPI_CLK_RESET_N
  PIN THREAD_COUNT[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 134.680 200.000 135.280 ;
    END
  END THREAD_COUNT[0]
  PIN THREAD_COUNT[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 65.320 200.000 65.920 ;
    END
  END THREAD_COUNT[1]
  PIN THREAD_COUNT[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END THREAD_COUNT[2]
  PIN THREAD_COUNT[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 166.610 196.000 166.890 200.000 ;
    END
  END THREAD_COUNT[3]
  PIN m1_clk_local
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 178.570 196.000 178.850 200.000 ;
    END
  END m1_clk_local
  PIN one
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END one
  PIN zero
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.810 196.000 38.090 200.000 ;
    END
  END zero
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 2.830 10.640 194.120 187.920 ;
      LAYER met2 ;
        RECT 2.860 195.720 13.610 196.000 ;
        RECT 14.450 195.720 25.570 196.000 ;
        RECT 26.410 195.720 37.530 196.000 ;
        RECT 38.370 195.720 48.570 196.000 ;
        RECT 49.410 195.720 60.530 196.000 ;
        RECT 61.370 195.720 72.490 196.000 ;
        RECT 73.330 195.720 84.450 196.000 ;
        RECT 85.290 195.720 96.410 196.000 ;
        RECT 97.250 195.720 107.450 196.000 ;
        RECT 108.290 195.720 119.410 196.000 ;
        RECT 120.250 195.720 131.370 196.000 ;
        RECT 132.210 195.720 143.330 196.000 ;
        RECT 144.170 195.720 155.290 196.000 ;
        RECT 156.130 195.720 166.330 196.000 ;
        RECT 167.170 195.720 178.290 196.000 ;
        RECT 179.130 195.720 190.250 196.000 ;
        RECT 2.860 4.280 190.800 195.720 ;
        RECT 3.410 4.000 13.610 4.280 ;
        RECT 14.450 4.000 25.570 4.280 ;
        RECT 26.410 4.000 37.530 4.280 ;
        RECT 38.370 4.000 49.490 4.280 ;
        RECT 50.330 4.000 61.450 4.280 ;
        RECT 62.290 4.000 72.490 4.280 ;
        RECT 73.330 4.000 84.450 4.280 ;
        RECT 85.290 4.000 96.410 4.280 ;
        RECT 97.250 4.000 108.370 4.280 ;
        RECT 109.210 4.000 120.330 4.280 ;
        RECT 121.170 4.000 131.370 4.280 ;
        RECT 132.210 4.000 143.330 4.280 ;
        RECT 144.170 4.000 155.290 4.280 ;
        RECT 156.130 4.000 167.250 4.280 ;
        RECT 168.090 4.000 179.210 4.280 ;
        RECT 180.050 4.000 190.250 4.280 ;
      LAYER met3 ;
        RECT 4.400 194.120 196.000 194.985 ;
        RECT 4.000 187.360 196.000 194.120 ;
        RECT 4.000 185.960 195.600 187.360 ;
        RECT 4.000 177.840 196.000 185.960 ;
        RECT 4.400 176.440 196.000 177.840 ;
        RECT 4.000 169.680 196.000 176.440 ;
        RECT 4.000 168.280 195.600 169.680 ;
        RECT 4.000 161.520 196.000 168.280 ;
        RECT 4.400 160.120 196.000 161.520 ;
        RECT 4.000 153.360 196.000 160.120 ;
        RECT 4.000 151.960 195.600 153.360 ;
        RECT 4.000 143.840 196.000 151.960 ;
        RECT 4.400 142.440 196.000 143.840 ;
        RECT 4.000 135.680 196.000 142.440 ;
        RECT 4.000 134.280 195.600 135.680 ;
        RECT 4.000 126.160 196.000 134.280 ;
        RECT 4.400 124.760 196.000 126.160 ;
        RECT 4.000 118.000 196.000 124.760 ;
        RECT 4.000 116.600 195.600 118.000 ;
        RECT 4.000 108.480 196.000 116.600 ;
        RECT 4.400 107.080 196.000 108.480 ;
        RECT 4.000 100.320 196.000 107.080 ;
        RECT 4.000 98.920 195.600 100.320 ;
        RECT 4.000 90.800 196.000 98.920 ;
        RECT 4.400 89.400 196.000 90.800 ;
        RECT 4.000 82.640 196.000 89.400 ;
        RECT 4.000 81.240 195.600 82.640 ;
        RECT 4.000 74.480 196.000 81.240 ;
        RECT 4.400 73.080 196.000 74.480 ;
        RECT 4.000 66.320 196.000 73.080 ;
        RECT 4.000 64.920 195.600 66.320 ;
        RECT 4.000 56.800 196.000 64.920 ;
        RECT 4.400 55.400 196.000 56.800 ;
        RECT 4.000 48.640 196.000 55.400 ;
        RECT 4.000 47.240 195.600 48.640 ;
        RECT 4.000 39.120 196.000 47.240 ;
        RECT 4.400 37.720 196.000 39.120 ;
        RECT 4.000 30.960 196.000 37.720 ;
        RECT 4.000 29.560 195.600 30.960 ;
        RECT 4.000 21.440 196.000 29.560 ;
        RECT 4.400 20.040 196.000 21.440 ;
        RECT 4.000 13.280 196.000 20.040 ;
        RECT 4.000 11.880 195.600 13.280 ;
        RECT 4.000 10.715 196.000 11.880 ;
      LAYER met4 ;
        RECT 93.215 10.640 97.440 187.920 ;
        RECT 99.840 10.640 176.240 187.920 ;
  END
END decred_controller
END LIBRARY

