magic
tech sky130A
magscale 1 2
timestamp 1608015951
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 566 2048 38824 37584
<< metal2 >>
rect 1490 39200 1546 40000
rect 3882 39200 3938 40000
rect 6274 39200 6330 40000
rect 8666 39200 8722 40000
rect 11242 39200 11298 40000
rect 13634 39200 13690 40000
rect 16026 39200 16082 40000
rect 18602 39200 18658 40000
rect 20994 39200 21050 40000
rect 23386 39200 23442 40000
rect 25778 39200 25834 40000
rect 28354 39200 28410 40000
rect 30746 39200 30802 40000
rect 33138 39200 33194 40000
rect 35714 39200 35770 40000
rect 38106 39200 38162 40000
rect 570 0 626 800
rect 2962 0 3018 800
rect 5354 0 5410 800
rect 7746 0 7802 800
rect 10322 0 10378 800
rect 12714 0 12770 800
rect 15106 0 15162 800
rect 17498 0 17554 800
rect 20074 0 20130 800
rect 22466 0 22522 800
rect 24858 0 24914 800
rect 27434 0 27490 800
rect 29826 0 29882 800
rect 32218 0 32274 800
rect 34610 0 34666 800
rect 37186 0 37242 800
<< obsm2 >>
rect 572 39144 1434 39200
rect 1602 39144 3826 39200
rect 3994 39144 6218 39200
rect 6386 39144 8610 39200
rect 8778 39144 11186 39200
rect 11354 39144 13578 39200
rect 13746 39144 15970 39200
rect 16138 39144 18546 39200
rect 18714 39144 20938 39200
rect 21106 39144 23330 39200
rect 23498 39144 25722 39200
rect 25890 39144 28298 39200
rect 28466 39144 30690 39200
rect 30858 39144 33082 39200
rect 33250 39144 35658 39200
rect 35826 39144 38050 39200
rect 572 856 38162 39144
rect 682 800 2906 856
rect 3074 800 5298 856
rect 5466 800 7690 856
rect 7858 800 10266 856
rect 10434 800 12658 856
rect 12826 800 15050 856
rect 15218 800 17442 856
rect 17610 800 20018 856
rect 20186 800 22410 856
rect 22578 800 24802 856
rect 24970 800 27378 856
rect 27546 800 29770 856
rect 29938 800 32162 856
rect 32330 800 34554 856
rect 34722 800 37130 856
rect 37298 800 38162 856
<< metal3 >>
rect 39200 37272 40000 37392
rect 0 36728 800 36848
rect 39200 33736 40000 33856
rect 0 33192 800 33312
rect 39200 29928 40000 30048
rect 0 29656 800 29776
rect 39200 26392 40000 26512
rect 0 25848 800 25968
rect 39200 22856 40000 22976
rect 0 22312 800 22432
rect 39200 19048 40000 19168
rect 0 18776 800 18896
rect 39200 15512 40000 15632
rect 0 15240 800 15360
rect 39200 11976 40000 12096
rect 0 11432 800 11552
rect 39200 8440 40000 8560
rect 0 7896 800 8016
rect 39200 4632 40000 4752
rect 0 4360 800 4480
rect 39200 1096 40000 1216
<< obsm3 >>
rect 800 37472 39200 37569
rect 800 37192 39120 37472
rect 800 36928 39200 37192
rect 880 36648 39200 36928
rect 800 33936 39200 36648
rect 800 33656 39120 33936
rect 800 33392 39200 33656
rect 880 33112 39200 33392
rect 800 30128 39200 33112
rect 800 29856 39120 30128
rect 880 29848 39120 29856
rect 880 29576 39200 29848
rect 800 26592 39200 29576
rect 800 26312 39120 26592
rect 800 26048 39200 26312
rect 880 25768 39200 26048
rect 800 23056 39200 25768
rect 800 22776 39120 23056
rect 800 22512 39200 22776
rect 880 22232 39200 22512
rect 800 19248 39200 22232
rect 800 18976 39120 19248
rect 880 18968 39120 18976
rect 880 18696 39200 18968
rect 800 15712 39200 18696
rect 800 15440 39120 15712
rect 880 15432 39120 15440
rect 880 15160 39200 15432
rect 800 12176 39200 15160
rect 800 11896 39120 12176
rect 800 11632 39200 11896
rect 880 11352 39200 11632
rect 800 8640 39200 11352
rect 800 8360 39120 8640
rect 800 8096 39200 8360
rect 880 7816 39200 8096
rect 800 4832 39200 7816
rect 800 4560 39120 4832
rect 880 4552 39120 4560
rect 880 4280 39200 4552
rect 800 1296 39200 4280
rect 800 1123 39120 1296
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
<< obsm4 >>
rect 34928 2128 35453 37584
<< labels >>
rlabel metal3 s 0 15240 800 15360 6 CLK_LED
port 1 nsew default output
rlabel metal2 s 6274 39200 6330 40000 6 DATA_AVAILABLE
port 2 nsew default input
rlabel metal2 s 1490 39200 1546 40000 6 DATA_FROM_HASH[0]
port 3 nsew default input
rlabel metal3 s 0 29656 800 29776 6 DATA_FROM_HASH[1]
port 4 nsew default input
rlabel metal2 s 20994 39200 21050 40000 6 DATA_FROM_HASH[2]
port 5 nsew default input
rlabel metal2 s 22466 0 22522 800 6 DATA_FROM_HASH[3]
port 6 nsew default input
rlabel metal2 s 27434 0 27490 800 6 DATA_FROM_HASH[4]
port 7 nsew default input
rlabel metal2 s 16026 39200 16082 40000 6 DATA_FROM_HASH[5]
port 8 nsew default input
rlabel metal3 s 0 18776 800 18896 6 DATA_FROM_HASH[6]
port 9 nsew default input
rlabel metal2 s 38106 39200 38162 40000 6 DATA_FROM_HASH[7]
port 10 nsew default input
rlabel metal3 s 39200 22856 40000 22976 6 DATA_TO_HASH[0]
port 11 nsew default output
rlabel metal3 s 0 36728 800 36848 6 DATA_TO_HASH[1]
port 12 nsew default output
rlabel metal2 s 29826 0 29882 800 6 DATA_TO_HASH[2]
port 13 nsew default output
rlabel metal2 s 3882 39200 3938 40000 6 DATA_TO_HASH[3]
port 14 nsew default output
rlabel metal2 s 23386 39200 23442 40000 6 DATA_TO_HASH[4]
port 15 nsew default output
rlabel metal2 s 5354 0 5410 800 6 DATA_TO_HASH[5]
port 16 nsew default output
rlabel metal3 s 39200 4632 40000 4752 6 DATA_TO_HASH[6]
port 17 nsew default output
rlabel metal3 s 0 22312 800 22432 6 DATA_TO_HASH[7]
port 18 nsew default output
rlabel metal3 s 39200 11976 40000 12096 6 EXT_RESET_N_fromHost
port 19 nsew default input
rlabel metal3 s 39200 33736 40000 33856 6 EXT_RESET_N_toClient
port 20 nsew default output
rlabel metal3 s 39200 1096 40000 1216 6 HASH_ADDR[0]
port 21 nsew default output
rlabel metal2 s 8666 39200 8722 40000 6 HASH_ADDR[1]
port 22 nsew default output
rlabel metal3 s 0 7896 800 8016 6 HASH_ADDR[2]
port 23 nsew default output
rlabel metal2 s 37186 0 37242 800 6 HASH_ADDR[3]
port 24 nsew default output
rlabel metal2 s 18602 39200 18658 40000 6 HASH_ADDR[4]
port 25 nsew default output
rlabel metal2 s 12714 0 12770 800 6 HASH_ADDR[5]
port 26 nsew default output
rlabel metal2 s 13634 39200 13690 40000 6 HASH_EN
port 27 nsew default output
rlabel metal2 s 34610 0 34666 800 6 HASH_LED
port 28 nsew default output
rlabel metal2 s 35714 39200 35770 40000 6 ID_fromClient
port 29 nsew default input
rlabel metal3 s 0 33192 800 33312 6 ID_toHost
port 30 nsew default output
rlabel metal2 s 17498 0 17554 800 6 IRQ_OUT_fromClient
port 31 nsew default input
rlabel metal3 s 39200 26392 40000 26512 6 IRQ_OUT_toHost
port 32 nsew default output
rlabel metal3 s 0 4360 800 4480 6 M1_CLK_IN
port 33 nsew default input
rlabel metal3 s 39200 37272 40000 37392 6 M1_CLK_SELECT
port 34 nsew default input
rlabel metal3 s 39200 8440 40000 8560 6 MACRO_RD_SELECT
port 35 nsew default output
rlabel metal2 s 10322 0 10378 800 6 MACRO_WR_SELECT
port 36 nsew default output
rlabel metal2 s 7746 0 7802 800 6 MISO_fromClient
port 37 nsew default input
rlabel metal2 s 32218 0 32274 800 6 MISO_toHost
port 38 nsew default output
rlabel metal2 s 24858 0 24914 800 6 MOSI_fromHost
port 39 nsew default input
rlabel metal2 s 20074 0 20130 800 6 MOSI_toClient
port 40 nsew default output
rlabel metal2 s 15106 0 15162 800 6 PLL_INPUT
port 41 nsew default input
rlabel metal3 s 0 25848 800 25968 6 S1_CLK_IN
port 42 nsew default input
rlabel metal2 s 2962 0 3018 800 6 S1_CLK_SELECT
port 43 nsew default input
rlabel metal2 s 25778 39200 25834 40000 6 SCLK_fromHost
port 44 nsew default input
rlabel metal3 s 39200 19048 40000 19168 6 SCLK_toClient
port 45 nsew default output
rlabel metal3 s 0 11432 800 11552 6 SCSN_fromHost
port 46 nsew default input
rlabel metal2 s 11242 39200 11298 40000 6 SCSN_toClient
port 47 nsew default output
rlabel metal2 s 28354 39200 28410 40000 6 SPI_CLK_RESET_N
port 48 nsew default input
rlabel metal3 s 39200 29928 40000 30048 6 THREAD_COUNT[0]
port 49 nsew default input
rlabel metal3 s 39200 15512 40000 15632 6 THREAD_COUNT[1]
port 50 nsew default input
rlabel metal2 s 570 0 626 800 6 THREAD_COUNT[2]
port 51 nsew default input
rlabel metal2 s 30746 39200 30802 40000 6 THREAD_COUNT[3]
port 52 nsew default input
rlabel metal2 s 33138 39200 33194 40000 6 m1_clk_local
port 53 nsew default output
rlabel metal4 s 4208 2128 4528 37584 6 VPWR
port 54 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 VGND
port 55 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 40000 40000
string LEFview TRUE
<< end >>
