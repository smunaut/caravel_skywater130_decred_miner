VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO decred_controller
  CLASS BLOCK ;
  FOREIGN decred_controller ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN CLK_LED
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END CLK_LED
  PIN DATA_AVAILABLE
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.370 196.000 31.650 200.000 ;
    END
  END DATA_AVAILABLE
  PIN DATA_FROM_HASH[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 196.000 7.730 200.000 ;
    END
  END DATA_FROM_HASH[0]
  PIN DATA_FROM_HASH[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END DATA_FROM_HASH[1]
  PIN DATA_FROM_HASH[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.970 196.000 105.250 200.000 ;
    END
  END DATA_FROM_HASH[2]
  PIN DATA_FROM_HASH[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END DATA_FROM_HASH[3]
  PIN DATA_FROM_HASH[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END DATA_FROM_HASH[4]
  PIN DATA_FROM_HASH[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.130 196.000 80.410 200.000 ;
    END
  END DATA_FROM_HASH[5]
  PIN DATA_FROM_HASH[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END DATA_FROM_HASH[6]
  PIN DATA_FROM_HASH[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 190.530 196.000 190.810 200.000 ;
    END
  END DATA_FROM_HASH[7]
  PIN DATA_TO_HASH[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 114.280 200.000 114.880 ;
    END
  END DATA_TO_HASH[0]
  PIN DATA_TO_HASH[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END DATA_TO_HASH[1]
  PIN DATA_TO_HASH[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END DATA_TO_HASH[2]
  PIN DATA_TO_HASH[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.410 196.000 19.690 200.000 ;
    END
  END DATA_TO_HASH[3]
  PIN DATA_TO_HASH[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.930 196.000 117.210 200.000 ;
    END
  END DATA_TO_HASH[4]
  PIN DATA_TO_HASH[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END DATA_TO_HASH[5]
  PIN DATA_TO_HASH[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 23.160 200.000 23.760 ;
    END
  END DATA_TO_HASH[6]
  PIN DATA_TO_HASH[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END DATA_TO_HASH[7]
  PIN EXT_RESET_N_fromHost
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 59.880 200.000 60.480 ;
    END
  END EXT_RESET_N_fromHost
  PIN EXT_RESET_N_toClient
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 168.680 200.000 169.280 ;
    END
  END EXT_RESET_N_toClient
  PIN HASH_ADDR[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 5.480 200.000 6.080 ;
    END
  END HASH_ADDR[0]
  PIN HASH_ADDR[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 43.330 196.000 43.610 200.000 ;
    END
  END HASH_ADDR[1]
  PIN HASH_ADDR[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END HASH_ADDR[2]
  PIN HASH_ADDR[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END HASH_ADDR[3]
  PIN HASH_ADDR[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.010 196.000 93.290 200.000 ;
    END
  END HASH_ADDR[4]
  PIN HASH_ADDR[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END HASH_ADDR[5]
  PIN HASH_EN
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 68.170 196.000 68.450 200.000 ;
    END
  END HASH_EN
  PIN HASH_LED
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END HASH_LED
  PIN ID_fromClient
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 178.570 196.000 178.850 200.000 ;
    END
  END ID_fromClient
  PIN ID_toHost
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END ID_toHost
  PIN IRQ_OUT_fromClient
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END IRQ_OUT_fromClient
  PIN IRQ_OUT_toHost
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 131.960 200.000 132.560 ;
    END
  END IRQ_OUT_toHost
  PIN M1_CLK_IN
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END M1_CLK_IN
  PIN M1_CLK_SELECT
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 186.360 200.000 186.960 ;
    END
  END M1_CLK_SELECT
  PIN MACRO_RD_SELECT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 42.200 200.000 42.800 ;
    END
  END MACRO_RD_SELECT
  PIN MACRO_WR_SELECT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END MACRO_WR_SELECT
  PIN MISO_fromClient
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END MISO_fromClient
  PIN MISO_toHost
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END MISO_toHost
  PIN MOSI_fromHost
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END MOSI_fromHost
  PIN MOSI_toClient
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END MOSI_toClient
  PIN PLL_INPUT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END PLL_INPUT
  PIN S1_CLK_IN
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END S1_CLK_IN
  PIN S1_CLK_SELECT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END S1_CLK_SELECT
  PIN SCLK_fromHost
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 128.890 196.000 129.170 200.000 ;
    END
  END SCLK_fromHost
  PIN SCLK_toClient
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 95.240 200.000 95.840 ;
    END
  END SCLK_toClient
  PIN SCSN_fromHost
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END SCSN_fromHost
  PIN SCSN_toClient
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 56.210 196.000 56.490 200.000 ;
    END
  END SCSN_toClient
  PIN SPI_CLK_RESET_N
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 141.770 196.000 142.050 200.000 ;
    END
  END SPI_CLK_RESET_N
  PIN THREAD_COUNT[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 149.640 200.000 150.240 ;
    END
  END THREAD_COUNT[0]
  PIN THREAD_COUNT[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 77.560 200.000 78.160 ;
    END
  END THREAD_COUNT[1]
  PIN THREAD_COUNT[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END THREAD_COUNT[2]
  PIN THREAD_COUNT[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 153.730 196.000 154.010 200.000 ;
    END
  END THREAD_COUNT[3]
  PIN m1_clk_local
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 165.690 196.000 165.970 200.000 ;
    END
  END m1_clk_local
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 2.830 10.240 194.120 187.920 ;
      LAYER met2 ;
        RECT 2.860 195.720 7.170 196.000 ;
        RECT 8.010 195.720 19.130 196.000 ;
        RECT 19.970 195.720 31.090 196.000 ;
        RECT 31.930 195.720 43.050 196.000 ;
        RECT 43.890 195.720 55.930 196.000 ;
        RECT 56.770 195.720 67.890 196.000 ;
        RECT 68.730 195.720 79.850 196.000 ;
        RECT 80.690 195.720 92.730 196.000 ;
        RECT 93.570 195.720 104.690 196.000 ;
        RECT 105.530 195.720 116.650 196.000 ;
        RECT 117.490 195.720 128.610 196.000 ;
        RECT 129.450 195.720 141.490 196.000 ;
        RECT 142.330 195.720 153.450 196.000 ;
        RECT 154.290 195.720 165.410 196.000 ;
        RECT 166.250 195.720 178.290 196.000 ;
        RECT 179.130 195.720 190.250 196.000 ;
        RECT 2.860 4.280 190.810 195.720 ;
        RECT 3.410 4.000 14.530 4.280 ;
        RECT 15.370 4.000 26.490 4.280 ;
        RECT 27.330 4.000 38.450 4.280 ;
        RECT 39.290 4.000 51.330 4.280 ;
        RECT 52.170 4.000 63.290 4.280 ;
        RECT 64.130 4.000 75.250 4.280 ;
        RECT 76.090 4.000 87.210 4.280 ;
        RECT 88.050 4.000 100.090 4.280 ;
        RECT 100.930 4.000 112.050 4.280 ;
        RECT 112.890 4.000 124.010 4.280 ;
        RECT 124.850 4.000 136.890 4.280 ;
        RECT 137.730 4.000 148.850 4.280 ;
        RECT 149.690 4.000 160.810 4.280 ;
        RECT 161.650 4.000 172.770 4.280 ;
        RECT 173.610 4.000 185.650 4.280 ;
        RECT 186.490 4.000 190.810 4.280 ;
      LAYER met3 ;
        RECT 4.000 187.360 196.000 187.845 ;
        RECT 4.000 185.960 195.600 187.360 ;
        RECT 4.000 184.640 196.000 185.960 ;
        RECT 4.400 183.240 196.000 184.640 ;
        RECT 4.000 169.680 196.000 183.240 ;
        RECT 4.000 168.280 195.600 169.680 ;
        RECT 4.000 166.960 196.000 168.280 ;
        RECT 4.400 165.560 196.000 166.960 ;
        RECT 4.000 150.640 196.000 165.560 ;
        RECT 4.000 149.280 195.600 150.640 ;
        RECT 4.400 149.240 195.600 149.280 ;
        RECT 4.400 147.880 196.000 149.240 ;
        RECT 4.000 132.960 196.000 147.880 ;
        RECT 4.000 131.560 195.600 132.960 ;
        RECT 4.000 130.240 196.000 131.560 ;
        RECT 4.400 128.840 196.000 130.240 ;
        RECT 4.000 115.280 196.000 128.840 ;
        RECT 4.000 113.880 195.600 115.280 ;
        RECT 4.000 112.560 196.000 113.880 ;
        RECT 4.400 111.160 196.000 112.560 ;
        RECT 4.000 96.240 196.000 111.160 ;
        RECT 4.000 94.880 195.600 96.240 ;
        RECT 4.400 94.840 195.600 94.880 ;
        RECT 4.400 93.480 196.000 94.840 ;
        RECT 4.000 78.560 196.000 93.480 ;
        RECT 4.000 77.200 195.600 78.560 ;
        RECT 4.400 77.160 195.600 77.200 ;
        RECT 4.400 75.800 196.000 77.160 ;
        RECT 4.000 60.880 196.000 75.800 ;
        RECT 4.000 59.480 195.600 60.880 ;
        RECT 4.000 58.160 196.000 59.480 ;
        RECT 4.400 56.760 196.000 58.160 ;
        RECT 4.000 43.200 196.000 56.760 ;
        RECT 4.000 41.800 195.600 43.200 ;
        RECT 4.000 40.480 196.000 41.800 ;
        RECT 4.400 39.080 196.000 40.480 ;
        RECT 4.000 24.160 196.000 39.080 ;
        RECT 4.000 22.800 195.600 24.160 ;
        RECT 4.400 22.760 195.600 22.800 ;
        RECT 4.400 21.400 196.000 22.760 ;
        RECT 4.000 6.480 196.000 21.400 ;
        RECT 4.000 5.615 195.600 6.480 ;
      LAYER met4 ;
        RECT 174.640 10.640 177.265 187.920 ;
  END
END decred_controller
END LIBRARY

