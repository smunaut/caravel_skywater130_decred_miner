magic
tech sky130A
magscale 1 2
timestamp 1608041000
<< obsli1 >>
rect 1104 2159 558808 677841
<< obsm1 >>
rect 566 2128 559438 677872
<< metal2 >>
rect 4250 679200 4306 680000
rect 96802 679200 96858 680000
rect 189354 679200 189410 680000
rect 281906 679200 281962 680000
rect 374458 679200 374514 680000
rect 467010 679200 467066 680000
rect 559378 679200 559434 680000
rect 570 0 626 800
rect 92938 0 92994 800
rect 185490 0 185546 800
rect 278042 0 278098 800
rect 370594 0 370650 800
rect 463146 0 463202 800
rect 555698 0 555754 800
<< obsm2 >>
rect 572 679144 4194 679200
rect 4362 679144 96746 679200
rect 96914 679144 189298 679200
rect 189466 679144 281850 679200
rect 282018 679144 374402 679200
rect 374570 679144 466954 679200
rect 467122 679144 559322 679200
rect 572 856 559432 679144
rect 682 800 92882 856
rect 93050 800 185434 856
rect 185602 800 277986 856
rect 278154 800 370538 856
rect 370706 800 463090 856
rect 463258 800 555642 856
rect 555810 800 559432 856
<< metal3 >>
rect 0 547816 800 547936
rect 559200 542376 560000 542496
rect 0 411000 800 411120
rect 559200 405560 560000 405680
rect 0 274184 800 274304
rect 559200 268744 560000 268864
rect 0 137368 800 137488
rect 559200 131928 560000 132048
<< obsm3 >>
rect 800 548016 559200 677857
rect 880 547736 559200 548016
rect 800 542576 559200 547736
rect 800 542296 559120 542576
rect 800 411200 559200 542296
rect 880 410920 559200 411200
rect 800 405760 559200 410920
rect 800 405480 559120 405760
rect 800 274384 559200 405480
rect 880 274104 559200 274384
rect 800 268944 559200 274104
rect 800 268664 559120 268944
rect 800 137568 559200 268664
rect 880 137288 559200 137568
rect 800 132128 559200 137288
rect 800 131848 559120 132128
rect 800 2143 559200 131848
<< metal4 >>
rect 65648 2128 65968 7248
rect 81008 2128 81328 7248
<< obsm4 >>
rect 4208 7328 557488 677872
rect 4208 2128 65568 7328
rect 66048 2128 80928 7328
rect 81408 2128 557488 7328
<< obsm5 >>
rect 226436 101260 229148 101580
<< labels >>
rlabel metal3 s 0 274184 800 274304 6 CLK_LED
port 1 nsew default output
rlabel metal2 s 555698 0 555754 800 6 EXT_RESET_N_fromHost
port 2 nsew default input
rlabel metal2 s 92938 0 92994 800 6 EXT_RESET_N_toClient
port 3 nsew default output
rlabel metal2 s 570 0 626 800 6 HASH_LED
port 4 nsew default output
rlabel metal3 s 0 547816 800 547936 6 ID_fromClient
port 5 nsew default input
rlabel metal3 s 559200 405560 560000 405680 6 ID_toHost
port 6 nsew default output
rlabel metal2 s 559378 679200 559434 680000 6 IRQ_OUT_fromClient
port 7 nsew default input
rlabel metal2 s 278042 0 278098 800 6 IRQ_OUT_toHost
port 8 nsew default output
rlabel metal2 s 370594 0 370650 800 6 M1_CLK_IN
port 9 nsew default input
rlabel metal2 s 281906 679200 281962 680000 6 M1_CLK_SELECT
port 10 nsew default input
rlabel metal3 s 559200 131928 560000 132048 6 MISO_fromClient
port 11 nsew default input
rlabel metal3 s 0 137368 800 137488 6 MISO_toHost
port 12 nsew default output
rlabel metal2 s 467010 679200 467066 680000 6 MOSI_fromHost
port 13 nsew default input
rlabel metal3 s 559200 542376 560000 542496 6 MOSI_toClient
port 14 nsew default output
rlabel metal2 s 374458 679200 374514 680000 6 PLL_INPUT
port 15 nsew default input
rlabel metal2 s 185490 0 185546 800 6 S1_CLK_IN
port 16 nsew default input
rlabel metal2 s 4250 679200 4306 680000 6 S1_CLK_SELECT
port 17 nsew default input
rlabel metal2 s 189354 679200 189410 680000 6 SCLK_fromHost
port 18 nsew default input
rlabel metal3 s 0 411000 800 411120 6 SCLK_toClient
port 19 nsew default output
rlabel metal2 s 463146 0 463202 800 6 SCSN_fromHost
port 20 nsew default input
rlabel metal2 s 96802 679200 96858 680000 6 SCSN_toClient
port 21 nsew default output
rlabel metal3 s 559200 268744 560000 268864 6 SPI_CLK_RESET_N
port 22 nsew default input
rlabel metal4 s 65648 2128 65968 7248 6 VPWR
port 23 nsew power input
rlabel metal4 s 81008 2128 81328 7248 6 VGND
port 24 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 560000 680000
string LEFview TRUE
<< end >>
